XlxV64EB    56c2    1340eT� q�#�X,b���/ʭR+$3Jçxh�������٩��׬}<%F��9�H�d���f��2�Я�E\o
x���c��I��E1�H�3��a��w�
:�u�!9QS7��
e���� �:����/��P��6�a!asL�e���V��3������O�NǠu��^,H���o�@�7��RZ�a}"Dr^�T`��8�*<~G5q��J2�K�,Є���������:\|R$t7y6�N���b�R�d%����$�V7,��R�ENX|�>εs�RE�l�B���5?�5)�~�c*4֐�^�@��n�1��s2>�lZ�&����B�.�e�m\ƹX�#YG�K.aq� ��uM�7R���(��
($y
��Oe�#����%HF�<�EC��%?"ƋK��,�%&u��?�=)�hUC�c�*�j�&b �Zp�O���"��T�@ޔ�w)`mVp����d�^�Ϸ��k�5U��+ُ��Voo�kNcQ�D�}�??��s���kLQ�Jm�Z�wT0&��{C����mb;��Q%R�Z���>#�$�	�CuG�.�z���G+�;��v�2gJ�Dh��r���2�� 䤦C�b*t�hD�M=Q���@���P�_ ���j̠Y��}�6]�rW�OdLP�
��!Z*��BA0����0s&�F���
$ �N�trJ�l��I��&�)��n��.�Q@l`ŧq԰K���2�k|:1(�F���o$;�vը�8�k�@>�Q�0Ž��M������R~RY�ܪf�+�E�%�r�y��g���5s��H���Dh�������e5�b$ �ܴ�l���\�S#B.O�R���F�"z�>�'���E뻈qs5��+G_�v9z�6������p����@Ÿ��zF���"�Ð�嵒{m�;��H��Ă����Q��g17�W�@���aɅspM�N�ԡ |�>I��S_�����5���X)�@jN�CX�Ө������T�ʡ�*��1QU��~g*zLY��vww|�M�(����)EI̭�E�\�m2����rR�8O��s�+�տ1}��g�0R�>q;��0�����)B��얳��4�ͽ{�*���4���cݠ���'#���W������w
���?B���d{��J{!��=�Y>�.�3��g��m���p��~I4����u�>7Ӱ8���sk�*v^IK�F����Q%�������mV�=�L���m�!M�b��nY��%�1�/ň`�8"�@�:����2�?��,�ó��ׂ|�f �CFC-�G��p���Rt��w���e-'�wN(�&I��A�����?��|�B���d� ���-���^,f���9�v��8�ǣ�Ŏ��� ���Q�zT�ʁD���5�ѝ�'��>by�]{/�
u���d�NqK��OM �^&jt"�B�õc�S��."�@�=�m`��:["���wݤ����eL3I%����
�q(-���o�庙)Y7Q3��]t�Qپ�a�&�!D ��Gev�Ɓ�\�L��(^�g�\�,MRcWP 4p�5;O�q�ݑ��L�³T���W.:��B_�h]���V�}o ds�� ��WaJs��O���_���O?0���B��~f��Q�IDȈO���y����,��'����%��jk��d��r@%[9��ue1�D֭ ��Qg�E�-iq�2I��_�����x.��n��u�P�l+��5g�&��z�z=�8
�-�$å%4�	�Or���"\��#� n,�tO��To�-[j͍g}lD��wS���8�h��h��R�n.X3I�_��7��ׇ�-��äof�����ib��&�!��c`�i|�u��$��=~/�l�	B8�y�i΄��`��Iʦ��1%��k�D��O�Z�DR����ŕ)6�u�:r���>�l����'	F+�Y�8{��|#�[=8_W�|E{DW��TlF;�I��k��V�*P��0d���m���M;�t��:&���U���>+�*Bt(򊩔46g}�����^��b&"���-#�eܯ�\��Yh$O:vW5��<D�^9+2TsGT�$�Ⱀ��C�g�j2��0%��Ԓ�IT'�j�4Y�oh�:��W��>�:���9�p�Qg~jD�W�F��p�Z:�b����i\�s�N��������v��M�xh�TfV`
��j�z���%q�N};��2�^�
(xzt=��}����@RWw�zp���Ǟgy�5�����mL�/JS�s�Í�� ����ט��b�֎�0��7*��qA�e�e�{,	�J�n�\���TAj�mH�}�k�"Gi0w���䂖�;�.�#�+����P���iz����'�;��؆�Ĉ(c�a9݊�Z��zdR��Y��ތN���+ i����C�誇�~��a%�ݸ�#5v�}������̱w���fRRd���I?��7i�w�)g2,<�m;�`�X
X4֦��R̊d�rmmQ�g﫢�������&1^�wlpC����~�P�Gz���~ݴWL:�w��`�"ɵ��Y~�����7X���7фOU�O��������,\gZ~E���թt�Gʀ�~���o0�fɝt|MY��_U��S�� Ȁ�^����_Z{�Y��.'��1����jc��{n&��C4N���N7}]��Z��Q�m��;�WҀo[YEf����s�u$;Oh����2�;A6�ŧ�J]�ɓS��=U/iZ�vǙ+?�H��~��"'a��y���Kr��:��K���p�Y5�Rp��J��>V	M�`�uW�[{�'8~��.(w~��u��Y0/G�[��LИc �?�0���j�	�u�kx_c�ʙ��͜d�0��"k���I�?n�����4w,(��6%}�ɪ����H�OA��}������i-�R�&<�1vx}ҧ��-��	�>`�x��	`��������ӫ$ Y��	"�6>��� Mo��å����)�tIA�!��zL��s`u9u�h��`�!P�I�.��E{�̧Z�\�V_Ff]�5�b�(R�#�K� =�.*�۾ �����
��M���ŧJ%N�/"���&v�5�Q�-�e*敵���<���C(�s2,"��̱��
�P��s�� :ϱq#��G�_`����kƖ_�*�����@#@���2��ʪ��@y{)���Xh�ݎ���H��Ͼ�,>��9�z�X�z��B��I�?¬xך��kɷ�s�5����}��"C��o�i����1�����4�݀�Dd�y�5����v2�����v�2��I!?���&�p�_���n������jķ�����q�g�q�ߊ�\; 8���$�Q`r(T�g�@bS��)m�}�=B�\jI��^B��ࠛ��T�'��3s9���:� 5�X�j��Q�OIJ%xL}�+���I-��RV��*��A+Ӧv.:Y��Z冾���)��c{�о����,�vUmkE��G�u�����r��=�ǲ�T6m.�[�,7a� �t't��������x��MBc��o����+!�]M���X���������'n[Qf��[���,])���֊ƺ���o���Rх�.A���lu^�	�W��V@�p��<蚻�{�֕U���]� 6�:AVo�saK��)kl�^�d���nA�j�R�g]��T��i��&Y&�b�d�t�R�vƋ��Ј��Xm�I��j�"Z������)d��cșBd�n8�81�)G�M�]��r+1D�@q�K��Ӊ�?�Zԑ��XIF "z�pL�JzG������+�g�"H\_XY>yݎF�4��=� ��q�C@Q�$H�&9a�zEUY�Y���6B�q�\�N��9�v|rAE�3-]�����`��K�!G3q�,�o�uA��_�	��������T�ܴ0;��̃��C��Ǔ#�f,0��ztXK� �r�ɠ��������u2����l�F<���੽9�MƧ,���vu��`(���Ȩ���s7���='G4"
����m�P��Z"�5�"��vv.�]�[�a�SR�}w���qj�4�8��x��sr�~X��y��z<�<�Q�>��qʰ7>�Ɖ�B5�#��=Yc hI�*UW�����9��s����\h�<@���`a?��5�{p���cu��>�4|�c���W��Kۀ����|�ؿw���ykK&#�dg���3�eT���2��q�q}���A_zf�V'�m(���ܲ׼��?A���)y��t�j2C��)��9�=p>O���W>�A�7_�h@�ѯ�Z�S�o��|kp�K�rOn1�����tu���#�e(���@������|� �w�T=o2?[!^{����/b�͞oƉ�n���3Y6 I�%�B ���9P�Vv !�8y�dA��a�-P�U���d��x���G]�X0�Ǆv��݅�,�0m^*I���B���,�<.��#o3/|�fgE!fA{��8g��a����	]z9�9��߳�i�-f��>V(Tĕ�_�	�;ǃ�,J�}ϣ^�qŇD�!� ���*��f�lif.�u�,84N� �нJ�W��O%QN,��J����*�l�=�{��$�׍ �X�D��H�0��{�3܈��~�	���-e�h���+�С$)���:Ѝ�
=�
̺y�K"��4���R�����Ҹ3���� ��K�����0#.qNe$N���`�U{��'DJ=]��@��} 4��{PD��?�?�