XlxV64EB    237d     bc0��EX���Z�|\�!4˲u�K�dq�ԫ��%(3�J�R���~�u���m�_�j��P��Asڼ�$FP{��oI~0��aܨ�]�
�u)p�f,�U���~�y}"����I|;t��3��V~(7�D>;2����b�v�&�?B�)L�o�#G��X9d��b΄8����H�@��*Yٍp�u�#�T4�-|�O����g�/f3����!L`�9�੟X3XT?-`��}m���)��f�oI3aH㽛ܗ�z�pE�u�������X�6���ͽ]����w�f9Ej����D�]��	��8��|4
��V2����6��2A�w�&��g�[^�P�r�] 1����b�6w7�ҟ�~|S����n��ߦ͎���;S�<f����8�M�b��9�̊�lCȁ���E�����Q򢌰JaH�W�ެIľ��qۨ�����H�����fPPi_O��$釿O!jdr����_�7���b��+�Mw�Fq��݇`ȓ��0u���W�K�*���ΡBڑ��^��a�wG�����;�3(ෞ,}�\oQx�I���%��	�T ��?���ޜ�9|�,�K���)u��+�~8b�g����q�������R�^.�>����*֝A��i�ؤҮ#��t���v>/�x"�����"�f5<bVT��O2s�%�g\�E�Џ�1��-q�S���Tّtk�B�\�v�u�����t�����(<x�����i����V�4"�z�S��U�p�����/I��X�ҳ�`/at���la��k��=��p��vN�S�W�>=�X���b�''rq�uv�mQ�ͺvݔ�R���~:IV��o�}��)
E]�X���k(��u&��!e��V�����T�����v!��[?>��q������C]-�X��y;� ��$1DӾ2��p �H�U�� ��p�d�$�O��|����y
F��n��#5�q�!��*�!��.�)o���+��))���Qʷt�>Uټvؙ��ۡ �%�`��B]�K39QD��psb؜\R8����,h��ѝ�+��BY�;zx��RVܹz���"�{̇���O'�`�T}�}[vO�,�xb�.P%6���ōcb|���I�<N�h�)�Dh׿�h;�U�?JA�%�!��o"����
��8r���*|P�x"����O��۳8
����b��cۑ�@�{A�Su1jZ�U9�ks�r�lao#$����+��&��m��o���d�r;qLb���v������IzZ���.dh�O�Ҁ�,]3��,[B��@�E��9���o�T�Ϸu�8u�cYN_��	����H3U�`ӉI��!-��xͮ��C�th�R��y^����s��2�[��H�)���nF,��c�YN�h��� �eU�)�n�(���͓�rc̈́v�U�ͺ��+����uO�Y���+��vp6�UKd�R3�44fo�ĥ5R|�%G�"�3W='jAaW\1�8�5Ǘ�K�I?�e�;ka?1u�!Ɋoq�����m�W����@�lV�͖1�
#���ȕ\B|��b�Q��r7�fSH&�ɔtqD�F2��{��B:1�,S��f��vl��H̒����X�'�����;R_�/�����n�_�XNx���|���_aV����\�L��������h�-�]�G��� �i�2O��X��!@U++��HDg9�y|��w�� ԏ5����[ַ���bo��kXG���1����-d,��	[#&��h��,7�P�%�L���T��0�١{�Qaj��E�o���7f�,U_3��?8K�`�|�4��eZ�1��q��;u�Y�JZdv���YݣmC���U�g�?WJ��C������V泀�^Qec�u�����ɐ1��8�mg@�|�I&�TG��W�gF�|���H��O��E����T���ן����Hط���0�l�@ge3���;N򍺬DM�!y��43��ޓ���ڎ���e;�"���د\�#6�|�i�c�u9� G@hI$l
!w�lJ��w���I�f8� �P�����"�I(a����	�� 7ϊ�Vv7&2�3�l�4w��=>�#HW(m�Q�U�Fo���X�"�VD�0�ioC8��.���ـىY���[䥣y�S
�;}�%�_F������9�P��>���?@]y��6[\S<�@>y0E/�'�=@�o�6^eӉ��"�t�$�œ��?�4��,�|�,!ia��!f�@*��#L�cG"�.�uQ:do�+>�Quݐ\hގ8��oLE�k�dǞ�}>�0rO�"��L�w�51;f�ky�~��o������~��0gA�|����9C��@�?rn��ѝ���Yn����%5�A�3s�^�?a��tw�+���E�n��U�7!Z�����g:���4�;��^yT=7�OY��Ԓ�/F��{$|���}<�Ȃ͏U��+�KC�_.	X�=q�KU��&��\i.V�zi{�!)�֥D��/�3��w��@Mhk�;��G��Mז!p��{\*J���.��T��C��}����&���C�[5�Y!��|���}��a5W<^�]PI)�$�l?j�&�ܷ%:�Y�r ��t���G�$,�	g�ˊ;�� �ި�=D����/�sMp��Ƚ��D�XG��</&�ր�w�7�8\�&
��R�ugy}_mR�ហ�����<�gR{o��$义��vӵ:.�G�~�p�kGfM�z��������O���Dw���1�wb���pg�}���i��B������6�b��ʟ��c�1� �#Zo���#�f�aϦ
�:��=�Q���[���|\��c$5IQ(-�"�%Ț�%պ��gXV��Qr�[3��L�$��{`��V��,�n�[X�եLQI�#�����,��S���B�+�u� 