XlxV64EB    fa00    2f80�bqeH�YC�%����%ʆ0�:Tj)��m'=��2����6p�@�I)�i���RYݎޜ%�/��q"y4�^�k�v�?�����}�����ԁ���'�����;,U�ӌL����r��{�߳��N����ok ��j�_���yNZ�R��7�5������ʏN9ZbB��KQ���*w/v/yB����0J4K��/A�nuRR��5@��6-S�Z|d�".����gQ,��K!�y�;$*�M((���ݹ`0��4���YM�'h���K���6)�Єu;L������B�cv�k����RgTc� ǚ�Y‫�ӓC#�{8W�q�'�{��SP^n�b��m��D|�?�!�!Ϸ�kKq�A;xKղ�M橮��CR �wdB�_��xzJ�8��|
���~!��>���6a:���_N�R���W�oc�4U���(��&�����H�id}�$����ʾ^Hi���AE]��ba��C^? ��x+"�UE���#}���a�z�V5��v���%����6�r���ՀX�N�-D4R+I���Jk�+�m(�_� Q�Y]HWI�.�R�1Fc9�KR���ftF�n�Uwo)E�4�ː�"Oe�Z�}�����"�D�x������qٸ�N�՟w��4��I�e�-��䑉�q%ZI6�/V.�ma�f�<t�ꓰ�}j�-�tp���l���r�UF�Ж�KU���2�`]aI]��,����e� �"@>�B�Yh�dk��f�9��[���y���qG��?��
�S�(D��o�����c� �b�d�ޤU5�D�s�0'�=�J�܋B�-� \��C�)���1zh�/�,]ȗ���:����	�G�x@!G?����kr���-�ᜳ�~�9��ǡ*�}���vj� �/n�;�#���Z/�S�"���]�u�12o�@bE�RvV"�%���HJ%&���帒��[iU�f���g:�o|�ܐC2�[�����E��`�i/\�8�Е�2���Nz����s��	b�}��!=;��o�h5f�RX�J�1��|�����>��O���/#��>ƚŧ��3�B���n��t��S�a���u�����a��[�8EJ�6�S�փ��Ac"v	�Ҥ���p�SȎ�Ho�mA=Ye�&�����@�Y����~{���i�� ���+�����S/��h�s9��i|�ZV&��1�Ɇ@�D�-y�����I}��A��8v���r��\"�95a�����i/���tY���G�o��6S�:�1"IX�Qr�kw��?�{w#��[�t�஠�r�D�+�����cY�*,v���S��rT�<��$`%Om9��q�\ω��
E[eir�X*vst1P��'�^ *m���T�?������?95�%�"<�pUz ��I��B�r�"�=P��}���C�� � إx�zb��� �}m�u�81�ޚ��[���kO�G� ����dcמ�o��]U��1P�|��K]��R�$�R��F��f�iTYbT[tq�?B��n�Kɸߌ �м��D����gOu�A�������{�E5��MȢӞ��L��Kv���z��e5����m8X�1+'�[��?�����9�T�o�6jV�3��%쇑Rz$�ȓ�X���-��٨_'~ ��^m�@R��sN�2F3�A���).����Œ�D�+˟c%X^����aB�m���k~�cH	�":��k��U���RPM=�+&cZ�ܭ.#I?�d#�N��[gC�
vl���tS)8�w�'��xM+�{���>Ӻ�M;�ޜT	�b�5<)�ן��9���rl�V�/BB��ي
�! �=�Cf+����~'���!����x�Z8�]�_���\���x��-[t�R@\M�GO���^IY�g|��d�;=�}�^)H��V��fc�$���˕eD����oh���%L�Xf��ϒތՎ��mľ�`4��g���K,M�����=�,N)�Cefs��"�u�&��h���R̓�Ġ��9P��ź��!�r��RiA�Y��AS�[SRN���$��BlD�����.ƱZi��n��SZj"_�R��H�
]-cr���˾z��+����>S�������bR��8e3OfE�O,V��Z�Wf9y���ج�|�n�}j�}݃�㴜#QMJ>���>-�=4��v�a�Y�Q<��d�eC;�"�cM��D�d$� �c"	�D]�r֔�y��ro�>1������U��Zq3���gv?���_���)�kD�!mHCI��-���T~�9���N�2t
y��n-w79L ��E=t�~�\��b��Y���W��\:DP����@���U~�6����A<X��`��)s��)(��[I|��A�()�!9��L<�N��'O)�(t�����g5IH�Вn�e$�D�m|fGK��/:���4z1X��{% ���i�(���k���e��G�3vH��Ъh���Y���1���%*���17T�y�$��ce9G&��d2�ܚ*�^q!n�&��N�Rv�4�݁^ �9I�8cI-^�6���q���޾R )�[;����u�`��9�����7-�*5�A�1�e�$�b0�{����M �$��Ƽb.t2�= yT��>��1��|� �
��'�(ގ|�h�44}����XZ)u�1�����{�Q��}[*@�w�ɭ�,������B�����+%��sR�Mg{ȝ�mq�����	�AT�4����W3��Jz0g�ٵ�"Y4�O�?�/���������E�״�]��qjXy֤�h�:�s��vE}�����(0�Pn��Ȧe���\���2�E렲�e̓���,DdN!%e>��:��Ŵ:Q���ʳ+�!d@�BKf����W2.\�;d�}����v�DF�[OZ	'NO�-�Xl�(�l2?���o�G��餡��ר�쩏��[��R�>WP1���F�d?H��,�*-2NOZ�V�@���+��&�Wefi�Z�x֪yg8�@碩}q�aZB/����i�ƾ�� ���&�y��e����f�Rr��t���Kz��K������(*��xG����N���s5x��S\G�[���E_�)��kC�=�=�;t����}�r~����s]�-���~H�C�)�B����v"��_�ƽ�<�I��	t���)�Y^"#�q9�m��=0��ѷ���{�8��"�Aɐ���"�TD�xZZ���h���>�JJl����lt5��s�`�e�;iPx���X*��ܕ�@�vx3��	MK�rk���CdJ;��KlF��{������a~+Y����q[��B���˲��a���n5 ?���A��^A�_E���]ٓ{�����Eoj̩@L8�W�i(��D^�t�}��tv_��
M�w�=��"�G����*�g�}���XC{���I��������mp)݊TÒ�Ežx��T��G���
���l�[�pD ���TT�o��r����z����j�����n��W�]o';RA��k��֐�Ӵ�dn���^�X1��r'8:�'�$mFŐЈ2����u"x�;l�ؿlk/��|!�B~�([�����&b#w�T�7_b�����΀�N��&ӂ��ROY�hs� {P�O�&�eSk��zP�i@�����6�!�����I�F�"����6��R�%�()kN-�k��vi s�[���H��q��Jmsw)9\$o� S�fI%�; vRT���J���+��q�<��Li�h!غW��i�&�Y���V�o��g����F^Z�#��%_1iKvz������:�@*�k>͕_�c�cA*�G��t�[�7��X��k���W��yU�:��
�XIyYgm�Q�����6b!)=e�Z�
�X6�n4�E��Ң��w6SC�֠/GAt-��l�d�y�낭�g_ib@@�\�ö;��zQyJsv�m|�Z$ �'M`��`R�9[�n�-�U��;�qΉ�	�>:��ɍ_L��4ɻŌ��E.�s��-%�]�3d�Lں��BƂ��`��;01�gl����!��r�R��)��g�n]�r�j��1庛�,���V��b>�)��Un�p�����iw����Ln���9��I����4/.���G��$6`N����&s�wuE����� h��S6+�Gm�d�ξ'����Qj�x|�k�O]F���駥�a�Gv�sZ���/ɱ �:!Q$��*מ`�� ���3��3�oë:dI��{`1��&)�2:��f+҄U�jo?�����l�8�4R�a��B��������ͥ���t�.��uC��Sʱ�F;"�`U�=�H�gu_�Ճ~W�ȤJO�_)��S=���j2��r��`-�֛j�՞U���l����j�6�z �K���a@��	� ��آ�HzlQ:w&��2��m���FO��$��^��?-v��Y�v[d�����:�M���<��q�����c�C��=s���x����E�o7��M$���>	T!����j9)Jm�Ű��-�s�[	��|�ٲ�����yw��sb�'ݦ?��&�O;��y�C���[*����:�<�'> �/e��45(�\��-��6��*�T%�^���t��i���~�f��b�~d���N�0.݋+�Ji�$�ǔ	)�h�axʴ%�F���V����X=j����_;�H(
O��g.�t��q��Ng ���u���$�2uP,���2Z�b��
M@D�:���� ���3�S	�����zQ������
���5\�=�p�j��G�?�\L'�A�Q����Z=�4|R�c�F�o�����7)�q������&
��|ݪ��>�'U23/
�Cc�A"���\��zQ�!�G V ��q�9�<����+~ ����xd�P�
e*=tQq�c�" �Ǫs��<�qy�AXAafLYp�.pkP>�Yğ�B�{&��+Hz SΣO��X�U#�V��TQ�A��m�H�?��p�wN3𣽎b7R����<��d���2A�$�ߥ=���[�Vf�`T/5�����(v����h+[�N��v��X����YIl��ݢx�^n��ܡp�u�Z���8<\4=�l�;�z�8�f���w���p�)Ń;%jD]�.}V>x;���l��cf��#\�Fc��hS���'�vU��˺�6* #��[�X-���N��i
��d`�_`��7Bx-mSª7.Iʶ����5FV�@Í�M��T51b�=�������(��y��=�g���b�L뙧-�X) ��t����Iba��(���c0�5�*��~N����eݬH_���.�&x�$��ʻ�FeZ�sk
~�A/�W^�j��C\H
���=LaG.㏺J͑�|6@6uP
D����I��-h8���0��?R�*E�1�}�ַanRH9_�ZWvz��è][��rt�����ar1��{B�Yr��Y^��]`H�)	���Ud2���9l_0\�3�'}(�����aey�$A�'�����`o]yl�X|��3&���%���l3�T&}�� X�*�W�}׎�(�(.�	��]kT"��t�x�%l�P0�7m�nп���L�x�M�^WAZ�3�R����S>[�B�;�O)��0�L�s�!(�21KM��Kj�T�"pS��N��<&��w��ɟ[�K(��ߊG��V��Lea�����7Ъ��C1�-��l�s���t:/:Ɖ��;�>��m�3m���7W6n�Dsܺ|RJ?F5|�-l�G�F��#_fe�F=�x[+eЭyWQ`��T]*u$���'뙃�\�����s���(�_���2����Nd>zd�����#v�͙��*e�~p��4uLg`�G�y�D��c����j�,�׋?B~<ٯs�}q�>W��Td���q��w%y�eR�\";��v�oE{_�^�O�K �9����́^�g�A��.����w�0ra�������}2Ͻ��|�z*�.a��a ��#}ji�W>T��)�:���0�"��(�Th�ƙ5�'y��v@
��'`0��f���T�ݦk��Φ202lIT�(`?a,�Q*�;I1ٗ���"S�Jv7�[&
^_Qygj�7ǲ2W]�sc;�������C7[�"����1՘��m�Kش��!��I
<YoM��A��෺��p�?���>ڞ!�uD��}���E���mH��Y*9�+�8g�2�a�ɿG���'�7+W�I�[0��X9�Uֶfa��V��H���8�p�� �^��\�9�`����yBZ
7[�,������I��m?ށ6���t6��k������+6ţ�{t�e]��㯺�<���FB|�����J����"g��D��ͺO�����X�'^h���R��P|m��-z�J��Ey��t� �,�If�.n\*�)2��4���$��z.��	Aŭ!��!��QE� �d�3������Qۨ�p$8"�Aԫ`�^믑u���gS��U�g;&Y�d��v������t��&J�ZE9q�F���¥��o_f�`�lX���l,����@�^�b�g�B�)����o��Þ�B���o
��~��8u�+��0�]t|�s(�?� �Y�X��<e{���i��H+��E�0��g�m�{A�r�=鱝�s.Eh�͑U�&�6�A��癯�#vT �z����L[�W��1F�W���T�|5O���=Kw���&���:�������xw;@.C����x*�:I�Z)v�A��1��[*$N�,��}������u�~	�^���v��岮�f_!�-���|����C�&�L��]���Ar�Y.���A0�'c�-���Z �[# B�.
�m�٫۶
n����x#M15 �Vb�`��{ �	���wXTJ,Ȁm.�R��gӄ�B�۬��m�R����C6��{�x.�^QJ�9HW�p3��͒o�3Md��~�*!G�Wy��!F�����LOo̶��+��F�Y@���$~H�l��I>���F�NU�(�hx]�{_)։bsj"�l��2��#,)��Ҙ��TDk)_\����>� t���dO�(<�]Lt�XOx�S�9׃��e"%�=���i��{�Ml�]`P24A�hO"�8�L��/��CD����y�Q5��~!?ˡk��l_�9�C�fz���um���ge;A���ع����@9f��.ęפ����b�7�Z,�#�����\N��=?.MmvL�@�bECB@Do{c���ـ�$�S����m�7%��UH'7��Y�/��f���*�@\�N�z�zu�_ �~UM���x�>6B mn Z��<���{��(pcޕ��\d��?��~|��"�R
��bhQ#�<]x�(��F�tX)�%@<�K0�x�M�1��=Xȵ<, 	^�]����x����F�q�0��j�D�����$��F��/��`����3��C��u��Ko�>m�]�JQ�9�^5�z2�y�9U������f�����2��<M���b+�G:�pU��M(�Dd�~�H�`j��:jO�93��&������7bѥS4'	�Y�Jkq�Î�I^C��v��{;.
~��}=�s+ۈ���՜���w���&�V���Ǜ��M��v�Q�HNL�CWE��5oD�40�������*�\���K�!D��t��i�)�>3QJT�d�P��X	��i'���m���8�k���Bͺĉx:��r�XPƝ�_k���c�Gy�5u� ND��_��t��+P�3[��쿺^U�?�p�EJ�b�o��{��%�Tu/`�_�xm.«�S�O#�L����x~��{�XQ��5�)[񀘲��:�5�u�ș,R4�G�Ɔ���6��L��*.��~"l����'cun����]y6�?h�ljQ�	c��Z9	?�ɥ^V�d3�~�n�q�b<�d~f�VF� 4[���免0@��۩]������CE�a`[�8(��E��#[?�K|Y!�I����锝�f~�8�}೔TTVP��5J-.?�_��Ȧ�]�v�\�.�!
+�C�E8��@7?؍�.+n��W^XX��xۜv�8�#y�̴[�#�����"'�yϭ�]K�H$�M+�N7���F�[e&��#<*�@A�tz�x�t-�L/�{*����+t�ri����0nrF���6��-��7y��r����>@Z�M6� �9=b^�=6���1z�R�&�e���+*���`�yv)c%��N�F�,�N.I�ۥϔ<W̮zČ�� ్��8�P
H��%'�t�֜�CJM��<�ܡ)���.�(ꡗ�P�PF(�&w���D`G�����A˶.�阡�A%��u	M�]�CCFh�6Z?�Z�h �����%鏿�Eh9�<&�0��2������N_�������+��8��ѾUsl��؍�S�%��ۜA[RI|4??�ا�>zw���RVi�Zn*;K��z���+�$2qA8��2f�����L n�b'�^m�!�Ȇa�����V�D��|��j1*k�Qi�Hw?�(�f���J3�T)�5��a�B��`(\y��:0��k�uT�e1����u5�1��Fw�~�u/*�E�iu�;d��4�[m�z��6P�l(S"-P2rA�e�;�54&�z�T��T��!�w��AD���n���wP�3� ,�ѦD�ȯL�JeO����]�qx�1O�����9�Q��0U���u�%�8�!� ��F���:b��tr��`8!3ח���$�qv禅}���t}�P*�}��W/�b�t�n��o~-;����-s*�ԩ��.a*ގs�-于���w �=J�4��'�\����{�ҤT�)��g�I㬦;ț���ߍPƻ��裗���6ξ�@P����Eؽ��q�k'~<0!eA( N��:a���T��w��֝���������mA��F!C���vs��Sժd�,���z�r����m�o%���f	�#y���-��T4&����˳��Я�CԹ�n-�7cX{��R�
�0V^?j� ��E�RP�ì.;�/,ޥ�¸�o7��{��'�}�,��!.�BˉiⵇWf1<�j@�~��~�{_���et��`$�a��⾱�paq ���j�[����B�/2���Q�i��N�~*8*%����_HB���\��
0:?��|�����b7U����>O�%"�פ<�T�mcG��cttf��!�w�`x���J�rRL�^�YK-��H7�w
���w��cc�*mW��MH��s(�W�#M��a���(,��A�1�r�����fy�d�9�)�y]w%Z�`�C��������vc;�H9_�pş" �.M!���Gj�ơ��`�xб$����4l=eN0��MMr0����3=ubHegѶ/i
q06���������89C�4,Mv�u���|���M�l��"���s rÑĢy��j��Rx#��8��2����?��Ϻ8���o(�Ύ���,d�o��?[�ڷ/T0�_�(��f����ngB+ҽ�J��U��$��b�n#�����t"	��ā|��w2�M^���bv���M�^k
.�0E͔���O�?F�Έw�I���UOn4Qd��?Kؐh͑Adu
�ϊ�a`0�ZCOP�; ��4��a�9�P�c�2k�,�����<M��+��Ѿ�nˆ�a�5�@uq�T����=����X[Ā�d�0d+���	i�Op�k���K��vC����
I���F$��;(y _��2�Tط�5�.�pNd[�����\�#�<���dCL�.g?�a�jA�ՙ��+ɥ����1�Vs������hvZ-���Y'`��,3#\�g�lu�-�����ʴ.�=EfNˮ���*�O��k���I��D���\��32����=�yV� o��>�(��sZ��-�9��������@2H�YO}Yܡo}�m� gj�z�q[�V�A �V�����K�5Que ﰗ���0Q��J�6�Txwf[f%��?��*Ѵn��T&��2�h��g+X_f�h&3s�����*Z��m[$\��Ԓh�pW�F�q��6��? �*l#�/P�<�d���^s"�N�K���؃wH�+d��_�sW�RZ�P�m�j�W�iiV�p��iH]�N�m
#	B{^Ol>JEL�����Q���
���\��7�(/��Ah03���w'�9�7w�V�]���	���2�bR�a�Q�t��7�c�6����F���`�ړG���pt��Zs<�%��(7��q�Gu��ߕK0�X�p���nl��M���/HIA�LJN;R�H��nz��|�8�Q��Z����1F_Ztׁ��Ab��Pq��_i��NK��l>/j/q�8�G-���
�gZ�'��J7���V�L�U*7��OU�w�Ѻ	"m ��	3Q�)���\�\�-���� {��b)�(K2���iS�����Bz���H�{�=�Y�K*㒕=��g�n_���X�t�:�ˌ������K�?�jZ'�uϴP���y���}Q?��d����e��v��&j;�c�z��QV ^�w%�#�EC�"A�f��m��!on��T��߫���l�h�%��>�Pe(��C]�s��5�ŏc��G'>'v3�C*��$��e)P�p�&FM�&���=h� �p�B2�Y)�HQĊ�N����FL�t֒������&��K�r}��	E�L��]ly�S��]����M;Fi���n&���q��� ��l-)m�I�$�q�P\�vȦ���2�����@͔�/����k��.����K#>����l�V�Yn�_�
��0Mbw}��j�5��aMj�.�	�> .���흪��-�f����0���i�|E��H[�{9	�m�7��T��DɁ#B9��tS ���n�MY���'�HE�������m� /ɧ�ψK�A*k��O���^l?��ur�r�|\7#ZI�R���R�@Ά�;��� �6:�) ���ž�yr��J�WĤZzE����fz�U��B�#�=����]��k�C�X��nM�m��KT2����Ś�#F��{@��M�g��j3�1YQ�(x-_�<ML
�ez߻���فE3�~��b˝���y�2!�+u8\qm�Fs<3/�D��.]��I�ؘϦ���*�x���y�g��/�H�	3�ܙ1����e�� 1�6b%N��#@��	��3�|W h���@	fc�¤*�>�*�	j�q=e��i���C��W��I�m7ۡM*Iׂ�"�A�­B��PB��+NB?�3��}�L�̒hU�Y�^#~a2�����t����6`��tl;t�F�����7H0I-u&ڙ2Kw��J�G�[[ψ�//�������H	a����s'�ꁴ���O
�����wU��#�*�ˋIDJ1jM^69�ie'��s�z����10�{� �?�$�b�Z<r,O���dΓ#�c�9�1�>����b�����?n�QG_�R��/vTd�[�O!=/�����\����U�b����J��oQ,�rN[m�'���Yw�-�틶uj��Y��b�΀Bo��y]U|���Ӓ+4�f��%�~�C�ۆ�{5n�C��(��ȌNO�2J��C���R-'���2��;��sn�)JM���S6��F��.�����3�B���j8D�:�SQ&ڮ
9e	He�|��i�Ϸ8
�2N�[pe$��A�ߝ1nbW�	i��^���=&;�DP�G<TG��̠Z�d%��=��Y�Y�=��M����	���p4�Ӭ1S����@�L}�HNas�0K�����;�6��:��!�פXlxV64EB    fa00    2b00N����[k��!�H^ ��u?(�3������e�+�ұ���J-c�'i��0m�!���~�+d�ޯLayw������o�Y^��k�>�W;����mލ���If��`$a�'��0K�Yy�M�dƫ������	*8z��{��!�|�r���.?LȋIug�j�N���7E����ˉa�.���� 2\��Ib^_�㎻��Vi�,F����ֈ��V�a���䓾��G.�Y4���r;"�Bd����*U\��`��F��z�!��a!���S�H�	��r�ې����]5�P(,,F�A����3����^��C2��"Y�c�u�f���~+�ydr��	@I����Pw�hqn�/�*k�L�)�#R+d�R��y�^�|�[�	Ȝ�5����@�M�f'O�q�j�.����͒�TX������NG��&B){�V�U?�c��(����mo
�]��Z,���j0f��}�;��>dK�{R��q_�Hs9���{�_����#�ޙ��7p6�Z�$볾���L�|��>�`�dW�����w��[�X���X��[��7젺*���C���
9!���`{�V�}�}:�}H�	�w�S)�W�2S�+�\�Xͱ�n)��&t�x���T}���m��z��Y�{��u��W��fr�ʧp5[���]\�t�*�"違41
�mjj:X��A���L :̓aK�q�ͱ��e�l#����,1=�X�Q)�p-sͭ�	t�Q~�!Ѡ4�-_V���Q]��Ѡ�'����iՐA
��	�\��)`tH�j��S r����E,��R*8}�&������a��V�;i~��8�r�aŹ��+0�G]�?�^3��%稆qa둣����c^ /;u��^�;�z��K�%��JT㦖��4�����'U�m�nc��>h�j�ͮ�#ͮ�S�\��� �va�țD%���H?�E���Yιx#�X�T��� ����Cn�s,q��&bR�ְ�Z�'р�2HvZ�SK��Br5k/0���p
�ti�=9"���t �B#YT��]0d!�H��U�����KAo�uo�Σ�Z�qY<��:Lw�e*�-C�W�vʃ��@1���B�?�ʟ��eUwۧ�)^n`  9٢R8Y��q��k�d�sk@}�X���<i �����Jf�ӵ���J��� ��_2P�=����G7�u��.�u����b98�Wџ�I��{��n�@�g��P�>�F$�8���,�p����F؛�&��Cp/�+��UIe�>[�����#JY�}f�+�ɕ&��h�j��9���[./�6r,�d����
�#`�ĳ��d�@A "Xd���4B�9�'p� 6�(S2�V�{�tC�lF���{����1h-�;$1�:[�5��wk��|!0�L���R��vu�:(���F�z w���`G�|��߰4�g�8� F]|?������|Ŭd�G
�S{�����t��aA$�?�x�?Č�\/��FT��Q�I��B��	c3x�*�EgC6{�b�y���hp��z`�5�8�OaE�4%�#������@.AlZ|0�)��F"�t�ǌəW���+v�>�%�{��j���|Sr�EA�(S�,�;���g5���Oy�(���X��z2?����kL�"��>�{u��Dּ�\C�=�
�'��ܐ5��#	,��^���KX�7�q_]�a��e�ӓ~�`d�ϯ~���i�*��%��l��4�9�=y��K��>3�K��A�£^�_�T*b�^V��!�ek�i�䪭w��Ԅ糣���Ex��$M��?A� ��2�Ǹ��~(�ſ��۝�ޓw��~�{�ܙ� K�"D���S�*�*�k&{X1"�'��1�$�}�od-�SE<�"�Am��U��� ���d�+7��\���t'�s��QT�v9`<��(F!k�f���9_��{�qa�eF��,#D�� �6K��
�L�KY�ӣ˰}�qr`�p�^�-����ox�'�S�)qZ�L�\s`�{[��f�|B��<"��,�PE#w���Y<��Q�%?ƌ�_��?w�J<�P���ݜ��gu_�#�Т��s� ���wՐؓ�^�Ɏ�z��apo�Le?p �8�ѫiVm����R$-J?��pY���[Y	3*E)M�P��<������i�����1�i7������}�jbsA=�9IY��U4��đ���Z/yEB.á�MK�ޝh�/�{��#Qm�S���4��0p�~8�����*�0J �"��wHHθ]4U8�x5��K{ք��n7y����?�f�v3�WKc�0���A�5I?����im��֊��'�!
�t�f���YPeӘć��}|%��4�	�f�76�����0>rOAh���</��!��^�|q�P�vi2קQ�M�Vx��t,�}I�|㘿��/�Jٓ��>�/e�lm�{b�	����]�l�4Ofj�]%)&l�6#��HA�M��-���w�v0�N,�W���I����i��4Ǝ�#g�V���?}s�vI8yp�8�d-�%���Z<:�'�����F��WHV��V����j�O�!�JC�+����&��#d%j�V���8��}�����
4�@+iIEQ�w�+�����RA敳a�r0�s�)"�n�̟�S�Q���������I���_Ѡ�Ѓ�_ۢh�� �U9Dڏ���q�0z���uH�5������vd�撋J;-�ޖ���%����Ί�?^ɥ��p�ۚ�d6��5�S�=�Pd�@9t�+"�����^��#Z�4G�e�{��Ԇ��.�l/��&}]>�����[O(��%�JY�?�8?�q� ��.f�P�[5����	��{��·����`'0�L��(6��V_ۭO�yI{{Wh�� ��0��V��y��<$��Y'l�آ��!�c��Lb���_��.9l)2�!2���-#šK�"��������L�rf��	������Qk����Ja��Z��jB �a"a��L9P�d��R��Є;�>&(<<�,����w��̩� M�6���C��i{���۝�[�}lV�'�$�n�t�o�~�r|�|-!y�l	re���B�*l�C9�	I�>��#bYT��� �8z|����&�E�E�!5��rE+�(,�ᒘt���Ƒ���L�
��V�Yuk��տ`]������>38�B"����U�U��2B
H=��;"ITt՟
@���=�^��ޔ�J3|�dC<��N$�yt��*�,�)�i�^��QR����(�/��Y��Y�$(�`�C�*�� 1�#?�rsv�/�C�ϝ[�����'t��B��"٨���r�1��a0�LW���.y�U��~ݹ���>��K��WV�P	W�$��VΕ�[A���V�*}$�E a�k�G~ �Q��p�L%#��tC7�̜)��|��+w��<��E��q�����?�	�;=D^(r�&!Q�	��|;�O�c8�̔��9�I}��ë�I��~��@ݚ��#B�U!���*߁�j1h��Ҽ����e�r�Tc�׋b���/fn�Z���7�p�&/�T��}���c�Ԭ�9�$Jm�]�&��n��>�p�`���h�l�R�`Ȅ��cV��7y��Gq�qj�s;;�7sF�;"l�h�����MA���'��3��>���k���pʯ�B=�GA��~F5�kË���e;l���� �q�X�U�jC:��j=�h4?���{!����^�_�Q�:ߥ�
�����[�AisE�tS��&�d�r���t�`g��1/�C�0n�ђ�j�	鑀dzPp�?�.�9X�{2ttNJӿ)���S��!I,D��H����8xx���v�2_�(7�NK$
�~�D��AG=ޕ�,^V\��D����9��E�of]IÃ�@���'~�+������8�9e�@2:�'�,��lh�Z�?��ahp����h袥�5�A:������&'"
��.��|'@(D�@kR���X�;����,*�1z�Fb@7�/B:й&`�}��uenx}iY ���d�H[E}���;�V3?I���댺������+��7�d�ղ��`L[�p������yeG�?�Wy�*����fNXQ�dEfx;y��D��3"�U���K� �u����UҪ>"��*."� Ѷt7t��$>7�|��d�Q�&�3Q�2�~��H4�̉�z���ݧ�Y��o� �&3�ex��Jm���5rLq��S�������� Lt�K�f6���;�c��"|#"m�Ղ��K-"D�aӑ���f
؏	�-tΖ�5r}��W�/`8>�c��D!�ӓ>Gx�����}�� ��_�+"&oV���)X���Q���f?sR����O��qڼm�=w_��'@��t�aԲn,��	}�9���$�a'���Qt��>,8v��{k$xQ�.~Ą���Z���Nn�AI�8�F��k�Ϗhu�v�gŀ.�P;���V-���sp}�z�|��b��E�����g�&�E��X/�<a��/>��B��ܗ'�h�dޅ?�+������ _�0��s߱b���X<�& *$W�y�..�[��lXs?���N2m�B�0U�]�oZw�Z���M�����.*�n�e�;n�RdvP����]�0Һ�tP~�ˢG�L�$�c6�3WS҇w13�'ɫ4o^B�p���M��.n/���Y�%g(�.���'|?yn4��d�
��V��۷,}]@��,�kWy�"d��i�[<ю
P���gR/��#�q٢7��]�ƟX_��~v�MEn-��j,��J�u�h`��4��6t�B��J��I���a��N1��+}2��eC.�-^�hs�#r_���<#�67�j����޹`H�6�B,q9}�v�k:���RM͈y�Eu�c�P�n�)�q�H�x�*��u�c_Â���j����<��4�N���$�	D0�s��� \���Jv!��-���lR�nT��?�!��B�����Z�8���N���i�"zL"�T�Y���YN3��7��vӼ��u�L�%��z�%ѳ$͝�����URTy������4iUE'Gw�Q�S�o��AO�+<=�fW����{�'���;�S�h�01��c�o[嵃��h_"��<"�熓"S�O`�:�sP�T�R@��J�l|Q�#���٘�|��?�*�h0a2'�[>Ӵ����R&_��a�[u�
�(� F�g����R�<�H��F�O�S�'D�P��5�]4��p"�*��9-�*�>Z���I`�'�5;�w�qغ�!�݁pq�a��&ht����>�Md9��R�F�5���H6�*&����ۢ>�~���D�$�`ۢ���=1������h��-AWԾ�#�V^�>*z�Y�8�q��u������A��SUi{��������4 v"o����1Ue��� 
��«3��?�Q���l���0 �"�d����J��$\���,t��r%;�ȶ
���e���h�`l�w"��^/��o�ؤ���H�°����(���9]�`k��\���[M��g�K P�:����6h�!o+e)��W��
�$g���r����_z6�PR��F����ژ��*��R�[!�Ks��!2�=��
sA!T��Ϛ�*����O�� 0��J����_4N~�i��'�^��i@<���kTT Ph��\����V}/�kg��K���s�§�;�G�=PD�#�|��w���)�7�����+��K	V�1wi,&�<�c �uB`/�84aMH�;����V�,�-ޥt�čM��[����8��@h�� r_��e�չ�R�<AkBà�EV��U1��nFS���:�H;0�@>�P���"���H�Ϗ�Hc��:��m��%a��)�i�c�����+�)a8v��.nIKJ�~1�aD<��w�K���@%o�K�t>,��`s��4���
ɏ1F3TO[�$�!Y�<�H\��5�b�@���J��k���iS��Q�R#aǩhyv[{c�
���nw,$�}�
��ӄJ�O�C{�}���(�H��}����f���+:C5i��x갏�F6���;�ɝ���v���{��Nley:oJ���aLT�~�pX����+�JӚ�?�ǲ�P���}��P�����%d4����"��,fx�斘�H��(Mt�_u}�²h[���V�P{r��^�X%����(���$U5.��
�#�X��Pb��:d%%+��K[�!����
H\�G��a����wХ��q�=�,@���ůn������`����?T�ű�Б��Y,x1��}8���h/ڡk�P��<KI�e�er.� h�g e�at��("뮷Kjƞ���ݞz;؟8X-ݎ��Eq�B�9!S0�0)�uI1�8?:�J����Ee�@��5�v��l�+��{|��Z���[���tt[��N����TY�?)�EhuI�4&�A����0ۗ�a�<+�����i����ն�\��ev����V���R�W�%��Y�˚ �qN\�����2��|�n��qږ����D®9�q�:�]cE�!\�L>|	��7x��#o���g_!��䒷<w}�-���2��e��xM��:S�t�w�	�'��i��\]�NM[�?����!�u���UA�dA��XH_APn9E��;r�&�e �	a�s���~\a�D����I:�<�u(ne4�D�RȨ��� B��r��]<ΓV�τpK)��~��yq=����᫱��������ּ������������i:�@����Z�p�k�̻=�q a�+�%d@'bތ��#R��/�:���A��Φ�LaI,i3t��%�L��\�D��'���&�BضS���tM)Qp{]�T|Kō��\��.��N@ej;'�������#�DU�0S��Ը�8+K��Y�Ŵ�v$X[���z��r0�{Q�`�6���А�C���"���#Jp�e޷�����4ȧ�_�	���C�U���DO���3$���QK��4���L`Ld4N%S�!祥��}�:��
��X2dA�ޘ�>ՐP%�F����a��YT��3���G�]��n^����S�	�_�$�^�?.z�����@G!�2��k�P���T�k�>�,o-B���M�&�.K�\g�\�`|d)��$q"����b[/}�x!@4|�,�LHM'.X��>Jw�e����Ѝ,Ʋ�u��~�ny�|Y'��d
:4w�+A��Ř
�|`A}�f��!����f�y�N�w��	�u��N�'��$�Ȍ��TӼ1����Z��3�x�$�E: VQ�%�)��r���٣�"����'�{�u��~��	-���-Āٲs���iNu�(ﲡ��œ��u�D"��3����]H�8��V+���"��F�C�ҷ�*A5�\�ĘT&�Dw؅j�ܓ0<:r5�f����!�]hC�eּwps�����&�SfB�Zb�.����� �GD*��~�^^Pv��W��י������i�`0�w�����%xj���DT�՚P��E�d�E�&_��)�T�x�
h#r%�A�ܚ��R���ڬ���:(+t����;�n�ά�؊~���Z�n������v���
bNU��z�̂}+ro��C҈TU���H�z��ܿo�����v��cw��p ��ֆQA�p8C7�/:��J�X2=�����Wk�����"��@��'5d��ucT�X��a_���M�gyT`������21�K�k�J�2R����O;�g�fy ������͏LDW��L;���i�`�qH��9���Gm�Q��3Z�k���=(5X�|<��6V�u�~��'
��q�W�Z5'�&�Q<����t
��X�����n��QS�Nǵ�
���;K}�pM��>��Afȏ\��K��{������<���%�ҟ�U�?=r���)K{SY �S����d�אh�k3��EG	�]�V���z�������]�z����|S�\� ���H]�wH�>��@��'�����_S!�HIk��V33Oe�r@����%�x��x�VWRE�6��1,�h��(+
@���!��2��'��\���v���V��O��O��68��]�v=�d[RuV��V+� y��l-���ܖ�(g/�a�Z�Z��ª��Ű�Zm�
<<yd$V-���D-�xn+!�00Ӻɠ2 �K3R�2�����G�$Q	/%��!e1��AH�?0z� � ���@�L�-9��>.�y��/�x��RH'��^��:؎���,��B���86ߙ��Օ� �G%~]N|C;��0�,����Â�@)�K���,!q�J���^��%jM�RŊ�N
��ɢh�w&i����,�H�ЯA�T^G�r�}"�p|�|TJ���2H$�E(hmhxK;��:�u�{���ب�o���3�#l{(ݚ��!��'x�]r�`C��2����c�BN�?"ex@���W66W�p�	|����\�����̻������}K������'��[���eS�EW��uhv�R>�Ϯao0�+A�N�'M�]�&b2W���t�_�&/	�id��4.��Xw�
oS��Vj�*Θ�s�)(,ȇ4ȓL�YVD�A
Lbc�W\����ԭ.����@���m%r+M�I��S��Q����R�<|��r�Z�*����e��u*��� ���j�-:�&c��B��`q��y	vc�v�=L�j����L��@��|myb��5��$�y�%��{M-;��G'�`6`���3�iZkI�|U�RU4/�3ɇ��.�����C&�:������[%S�r�z��Mz2��"��9ֱ��g�K���OX���)�Oi1�g�83_
b����`�C�En�x�#gjϑA���#�@�ϳ=h��\ac�%(Ne�h_V�N�^���z�6�Ũȑޚ�Q~
!J�T��P��l�[��Ƞ98�~�2U����@? r��fSdV+��/პ�;��}=���8�n�"l�4�H�bkD #{�A�+P.����]b�=�ւ�4�j`�l��|�-�ޫ�dB��!((����Ԯ��^Z�r�	��;��Yb $αЯń
�	x��Σ�h�@x�H@]?�*��

_.�R�a6o�G��}�� Ow�wx_�}�ր�R�n�`���d�T����12ѼuC�z���n��J�7$|l�[�)BUv%ym��<�̮�%Q�����t60����v&@h�����{{M`C�		m���M���Qh�T�E��٠A��'��N_k+�"���5�x�J�d5�!��^pj��}���'��t`�T@Hw�J��T� 0��D�V�$#�����I��+�dc�r�����i�`�YR�|'l���4aY�ӵoe��r��]�F�eb�ٽ�2�uص��t��!�VW���I4�ʙ�o��c�����hFK<}���]�����TĐ��4(UT"g�:�%���� n~�Vǔ嚼.���N	����ZȐ�a����{L+FB�����۔��ѧ��('�-�N#|����_���LV�VCpV��z����{~�����Dݤ��P�t9 E]��	�fS��-г����������t5��V�^�)�w���A����y��F�Ys�ۋ<����������e��a��fQQQ��nS�q/�fUQ�H�z����1؆�u��]z��6̟[�t=x.peg�ä�&�7�aŻ6��}��-����]�5����Ѕ�G���&���U&��5�ărg�`�����Jk�Տr�6��r��C_��?�G�|��kPE}��+��ʃ6l�~�����`�酴�J��[D��K Xy-�\o����%�1^����!� ���G쇌[���zi���"|�[C&ZT����2�x��o�+�͞�����^�|얍�&K��S�꜡��C�D�H�܌�z�K��W�T�.��*佼�.2h�#7��dcp��_`N�,G}*3���v��"��ܲυz':�蹊!׉�|@#�G�v�ʞ��(l�\��Oyu�$�7tpB��:^�o�"~@D5g��rn�^���-�y܎�Bj~��s��j�`� �3��z����Hk�F�ϒc�0���`����c]ٌ�xʖ�$��*��vEP�nCu
��Η����{����{�Z/�p�ڱ
)�pVv�^�*
�!rm��Yt��;2�N'�B�b�x���Gb��"���������u��9�r��+��B*f�nl����`�f�-�G6�4�a��L����9���P���iJ����!����}4��㌀�k	���N�-���d8ԒE�u�c	z0��8 ��m�>p��WҎ,�j���t�jE!M��>�+������d����+��SOX��7�p�@�m>�+�PM��n�nD���Jy�g�� �K*��Mј�arJu%
x� ���5T�͞J��2cQ����x��sJ�n�@C�ZA����x}���O0��_W�p��Q.�U�qW;�1/��]����8���(����"�A����͙�VG��J�`��P�,t�TRv�m��fjy�t a��{Er���b�-ӏ���]<`�5b"���@R{�Z�8��+�Hs��2��g���'����O-�N�Z�s�4B����N��JR����z�E�Uv�*���[
MHv��8SI�7u��:��@�n�po��e�%W��=PlV7��*���& :�\���XS����p�	����ZA����0���3%)�J+�'R�;�Z���`��
hYe��7���!�2�����CyWò_Mk�_c�_Xhr�J��9���s�>�I���>_m�/}5�[O�XlxV64EB    fa00    25c0k5";s��"6f�7��G��^x�**�(�Gᛜ��`E̟�D�T��Z�U'�y)���-��mE�H��GXHx"��6���P�c@@&���v\�+��5#I1ͤ�L�LDHx��VU'd �U�Z�����B�e7�Z+���o
��F����G�af�'��3���Vi9��N���o�H��e]î�}�ӞtG/���~�j2�b4Ɲ0+Ja��ۻ��Ȭ9�H�DAĽ����`�`Ͳ����N��moR~1n�k���̌>��R��isv����G��>"���C|���\<%�O�#՝M�&rM�i�� ��ظԅ�g��O�2��m�}�ëꛐ��iɯ��~�Pt��/`��u�"y�n���O+�4�f^,6����Dqb����n��\��g$����2YC/�nK��4J%� ��k��9M<�-��V_�0��[�,��>�x���_���f���Fm~'=^8���Zn��"�f���*0�Sgߞ����fCJ����|���2ۼ8�9�x3�؞$
����, w��*�I�G�1�Z0a�x����Ph�'VQ}�^�I�tq�ھ��O��T<�"�԰�I�n�q�)^~�dZx���Kؙ�x>猠d�ʔ�2�%��զF��ڌȉD�Ph�B��� �S�gQ�(*�$�$]LK����i�t�܉ۄ*q>C�E~��u�^`����>��n���nT��ۥ�E��F,�	P��Z�']x{��^���g��-����'7@����o�8_E5{4"]DP�����Cr4A�&�o�O�iٸ=��1��F"S0��7�DvT��(��I�Y���8��|5�"\����|rM�9��UA?��3ꛡO7�m�/ -��.F�C�ؐ�Am�Β�${ݑ9���4������+zzf����X��V[w�#`	�A��c��̒�a,�3���y��r؟��V22\i ����m�?��y��0��;;�Bm��X�+���8h���`��c����_��h=*5�+;�AJ�:������#���KMR;�	�V����'�R�XXԃ�V^h.z�����AN#�>^�9`�̩W^E��$ڣ'vTⱣS?��Jg� ˼i�!s�1k%�[�5�
=I����e�V��:�C%A�	E�Xw����:�kHK��4�^q�0��[p0+ƕ�BH�]�<��߭�vq���HMk]2��"�Q����6$� ���SRV�K��[�a���*࿈v�*��=Pq�='�� `H��I�x����@Qɡ�G�=â&�wc'=eҎ��o�ً7�\D�b�Z3��K�i�`�-�����wv��@�UK��������AM�Ba�_�R�KtmM�[	��~K(7j�3)�L���T 3��\DE�;j;��DmX5_���r�5�HU�I�ʌd�l���\�9}PO$>��Q�M�΁ @� ��9�N�u���� $�A]�.�s��q:Q�jf���"� lq�^��6���"ԏ�q7ơ����kt,�{��V *J#جy"�%�8��A����|�~��%�5im��F��I�*��b�ݩF��-;��F�8p�tJ��׍���pU��>�v=Kࣃ���)���8�<���w������u���OO�����h�?��g�d[z��?�EK�ڹV��"�H+��S�X�S� Ml)������ �2Or#�ڌ����p�v�b-����|�y�P�lc�7�A_ƘZ껑ۼ��z�&�_�1e���ao�ʇ����S�9T����<��ѫ, x��DQ�@���|ʜVM����f�����Aϵ�8/��y�ZZA��s�ۉ=�������d�d3��O:�4
=�R�7(
@���_��Q�M��0�����y8,�6�T'���L,XjK���^��sY�hE�w��D*��67xw��JɗV���q���YD��}��3���D�]K4G�w���u%
��)��5MLUm�]J;��R�a���7l(�3�'��Ç/mH��V���cf�� ��m�5󔖸?���V�ۭ]�&�isJO�}��k����<�&j5�vF!J�M�p��%��نB�A�1��e�%Y��"-a/LЯ��~]��� y���������~�gD����ӖJ���^��t�
��Ұ/z�י�q�*S+*�O����㈸����g��t��T���>��<*���������0"jr�p�*�v��HyFe�Lp�J�"����+v�݁�έ��4�"ޛ�z�ևYvr�<Q����g�y��:�����[(S���4}g%� �}?�`���[[�(��O�77�)58v�w���ɷj9�O����\tW��?��e�@�&�M�J��'8�Tε��s��@����2�`ĸ4�ך�fÕ�m ����gZ_��� d$h�[���]����v�姰9�P�GB�.�Jad'�R6��L���9"h[]A�شÚ|{����Lh��F]��ޏ4�5Ry�����3K# e�����;׽�����`�,�v���ot�&4�,>;ek]fސ��٠�fm��Q���2���'��k�4�!v��߾PpL����Dm�<��u���ة�XU�+c�3��C���#�;��`:���W41�ݜ5%���<��39��F���,G(�}��U�o��h��pbh�4��"�į,{M�p�d�#�'�>~�`Iw�ɛ�)_�Z�,� ��C�7�t5��щ����g�`���>�8w���1�dP"AQ�Z��w�H?�m�	6}k�Z���Z�*c5�+��tDS��so�
c"m�GP���n�N�������&*R�
w���{���"����F`c>G��W �+��4]�O��X��[�77'�ğ�'���篨��������6a6Oq��K(xw�P��CÂ��c���	X���*��:H⑻�"�z�D��5�%�Z���:Q��h�v�h����g�|��+ضV?n5�:�ܲ�m���� K���9Lxe�Zb~b�U�}�n�p@�:��_��@�i��ˬ��A��@�4k�]����Ӏ}*ѵOz�Z���Ĕ�w���r�-D+ubY��#�k�! f*���{Q�%�74�}�]8�G���ƴE*�����>Z�K@�L>���h��=�V��?����������*[Ml����ǲ�8r�� }����iI6�}�u,ɐ2C�������,���>��3_�iI�g|`����u���s+JN����S�Wu����4X��wd�������@�,�IN�
���\��o�A�g��V�P����$S@��{Q~�0cު؍�Z��o^+��c�	m�����+{'����J��')�����Al�f���f	b%Qku�D����Dp�����r�e2��th�nַg�U۷}�N��k�� �y��=��f��U{_���h�AI��'(�9��j1�]b���Lnf��xP$Q�q��Tjq������g�k�
K�<BD������Gr´��ܝG�nl�������D�4L5ݟr�_�Y%�v_��<'���/�[�yH'ʓ�Q�5��9A������z����=�`���a�1T{w�As~Z���-B���H�j�O�x·�t�[8�a]��-ч Ȥ(��?C������:�uޢ�&�0��������!����w�����o���H2����/���b�?u�)jdo�������� ���=��?�C���@�#��\T����[[��c�O���8�x���; V��'�����r	�J�cgڷmh+�+0*����>���ν�+�9��g��9Wϯs�ڊS�d1LB�G�d������6,����U����UG�:��N��S�L	���L�8��؋`�nm���Kj����_
�I��`�}؎�֏�7��J���1��ɗ0����w���dbyի��Yd_f��ފ�����;�ϟkk���p��/5�"qJ��F������I�n(�؂����ؕF��I�����n�q���z�9 y�G�o��̣��^�tT[�o$)h�ьOǈ�C�L��������)W7!���&H�a�_M�o(�ط�2���*m���*%�h���I5[�ĳg������ ��n� ;i["�g�|��{�������f\��p���u�g����%��7j		����"�J���l�kܗ8_�<�k��������U�%r��Hˑ�2���!��`wb��p<��^<��J�x�6��t��'L3�*�>�B�u�(<��)��!.��W�O�>�#��{�~�O,xx���}�����_ ��J·]�43Ԟk��9��D�4��x�t�V�·�L�Y���J ]��,�;y�&,dua�u�iG�f��[��c�Gj]��/�	l$>�)��e*���\����HP�v����ܜp#�L��z��}枲���)�EXt��KI1]j�����n��i9��l�7��&��[ h|��U1�	Fre%�Cnx�r�h0b�I�$OE�y򅀚���+�hVB~L����e�$�/�z��ج8Ⱦ>vϊ���b��b*��)ד,"����î ����;}XrU���P,'ɬ/:�[�WG��:*BI��l��~Dj���Ǎ�`�Q�
��JUg̱����rVhb�u��h(�5`�5(�}������� ���%},�լѡ-�]�]E�>��}�uq��z;�ϗm�Z��[��.���ᥓ�==�oX�L�`��^���I��0L�Ԯ��`pӮM��E�*�G�k�z��ř_r_�59@�숋�U�&�q���5��/�ߛ�cJFS[��ͻ�)4-b�K!7Q@����X�������Rcw��f)��INP��JE�	(M:򫶊%���N��U٘�7C� X���܁�3d�B#K5�aߺ	n��[�OS�zed��#82gN�V�|�G!ȓư�z ��]�2�aT� B�Qf�<��oRw��2p���>���*z���\4�_Y�gֿ�
�~ʫCR;^q��`b0g��H�Z)>���F
�s���{ޠ�;o%��jT�5��"�Ǝ�������P��Y�c�l��9j�RMPV�>���'��a���J���/	LȽ4�����r�TE�֐��Y����`z&������4&)�N�y��%2�� ,T>��|J�e�a��gY�٩-�g�Mj&3G�ި��0sf�<�K���ʅ��������0wH/[Hz SʱԷT���œZoɱ00����.弑��:[�:@���~�u?MM^�)Z	.����Na$���\�-5YH(�H?ġ���cU��������Տ����0V�����"��T�3A���X�P��򜅑�
�Sσ�]�GM�7���ɵ5��<|7'%��A�IfW��b�b���Q!�x`/�"f�pA3�$�6�T�{���#�t��
^٢��d���t ������4i�⠉^�qP�Njy�%Ӭ���OPړũ���LYe��B�O����;���/V�� s!�(Ǚ�W���j���[�E�$�,k�C�^u%�b�G8fH/ dT�mL'^���lޖ|�E�,[M.b���S�|�T��񜵮u�ˎ_\)��5��=|g��9Gc}rp�Ҳ�;ڤnv�%�&�|\Pݡ��3z^vl��5G� ^�[b���ou�iqV���_�X����I�P��0���#�Y��@)��&�O\���k�zh��1�M��Bj֒�-G��^�E_FD����	��7��$���RN�U�X�g��@��=��#lĖ�{�,�7I�H�碽��K�..�L�FxC�6�HH<w��$T���iк���*I�bd)�T��1˻��i��g��a�8�j۽�v�c5����|��R�\���:C�:��z���vx�W�)�+���3�0�@�^�qL�����1M��3�$E����Т��Y�)ƣ�R��g�.�Qn_��p�������f��2UV�|5����o樓="��d����L��({{6��T�r%��ƫښ�Oʸ4��[�������i�_���\Bߤ�XgY��A�1�����!��׹����+-��:�Ŧ��;�E3�w��g-��^]K��Z�5#[��)��3�zd���9��+`Y�N�k�e/��Q���ҋ���9�������ݻJ�sq�~���J�uu <����	0)tK��'�)�y�:�N�P�̀9kTj�&�6n��}/*�o%�Yyb���yK����,��&bN�TЀ���#������s�/{5�D~�}V�B�,Q�Rּ��o�ջ��FT���Ak�V������Hz�"����2?�JQw�2AF^�� l������ Wq�Z��$�7 fg��?�!�P�׸�;i"{W�̓��9ܾ�D$��1˗�Ay��!�S A=��r��9�C�^K�@��15ޫa��ɛ�bd�,�.��k;��|@����&^Mx�2�0��&�8 �.�G��yt���p�`�fkM^�#�*Uy�q��=6JM���u�vV306��Óz4�[
���0�$�%S_\?b�pҁ;Wo�{i���+����4E9������vsq�+�h]@�e���aY9��_��G~� ��ل�;��Z��Ԋ��Ɵ_e��Za�w� pN���}�=x}Y�Ë���_.-�h?C8�D��	LR{a\���_��e_�� �X������	�<��p��hH�ov�P7�޻g}�/�
6O&2�gR�2,e�0�S`.�SU(f��\+��5���_�"G�`�X������� Tg���T}ך�L��i�&7c��׿�4�W���F��e�[l?�Ǩס�E\ ��Ux/����6�F8�)ѡ�,+��jQP�{�E	8�	`�pd��{n����a���Y���u�s���V���iV�^������A��"՛8��^-)�1��щaq�����k��;j��(u�����.��T�&M6�2��'g���,��LKc�V.z���?��Ŏ�f��]�N�x����*��2]���9���G��X�e�p�e�f��� ݧD����0%�Ψ%:�
m�+����&��]�
�_��P��;��� �9����EN�i , L��0��_��߈��0اx�^g}��d`ܴ�ǫr�@���*��p&��
���9�����Ǔ?�E��Z�X!��^C5�zF�#n�}�m�p��/J�8��q{��d������s��������ab�z��Q�6�`6�Je��O\�Ge_���g��7�����c��r����/qBZ����W^Zh�X��ξ60�,����}Ǹ�l	�v��z��W%˿%
�]O�G)G�㰮�\�t�%G��ЎT��������Xv_�R�
�K@f���ٻ8��x�`(�'�>�oO�QײȊ�S�������N��p�uמ�^1���+j�6,��);Y4��c؈��q��AM;��X��ቬ)S����Q[�R��Vs���*k����6ɖͯ2���~o��&8J��Q�@�z�$6�*ÐG�n#`�m��k�ܟ�Hf�s�����o��*�<F��ba
u�K�>�ĵs侊�-�0bK4����N����*�M���jzށ�I
a�;b[�_�3�X8��*c,B>Eٚ?H�2���8��%W�ا�1z�Y�>���H�j&��^|�2�n����kV�,�c[�-��0�����Z(\l���]��!��m)j�t/@Vו���0)R)�=���qx��_p|G2_�T�QY1�5����4g�湍fD��rI>���fb�� f�0»d�b�埱,�ń���Qɹ�m ad&�>��,��w��]L�J�����G E����iVfw���`��{*c�� �v�$����3�[�SEKe�A1YO����"�����X#�p�ø"�Z�͵�]'v%��VɽI�!B-����B�b��	qk�����g�eS&ơ)x�����-��T�K��I�H݊���l8�壀���%ͫ�������W��ЦB.��<�e'b�(��ɧ�������"���c�h���-�x1����y�˩T�3vI/c�����(\��i���*�-W�[\��H,�����B���E��׺4f5!�5��Ǜ��[�7�0�"
2�)�\�&,�;q��|	�r)ݶu��>���2��@���ދ-�pb�� U\B�4���vi��d[�V ?�Jw=~�BAJ�rs�b[:�rd�� �e*|z�C{5�x�S�a�a�4Ca�����.��靯fG�<I�+ce�O�����}��4i���K*�^k�X;��'�`��>���t�G\�o^��"`��֗ڞ�y^<�����[qfٔC�K�a�tD5��ө�A`H�h�6֐�Eo�ztᢱ�a��,a+�^!��K��kh�Td익�!���	�9\C�<�[��i&�������5@�&/���$K�8�cX�R	{�&�U{nd�I����*�<�b��b�����>/r����Z�r�9��X��L<�&Pw'�R�%�����W����&r ��K�d��� 5�� �Љ� YRQK�T��H��k.�!J�0���D��c�
�9�p�A8l�!�aq���a(��6_��lv;vu:��5H�:�2
D�Tr�t��&e��6�O,�t�o�p�:��#�%�<��J�3ۧ�sնW}�g�n�#F��S��P�ȯ�(��� +�cՕH����8�[Y<����{
�po���0#�[��O������
+q��흆l���#������kU���0��ݜYy�H(8A���:9�;���vY�Eҿ�sc���?;E�KNL͏	�P���H"�%8��TDE+r�H'k=\.nÆ΢ֽ�|�Eg�^s��Iw���X4��g�Y���z���l:⡑�M\͟wV��w��	O�G�(�F������{��$��F>.�cyo�GF�}g[m��Nҫ��.����8y&�,b���ƽ�{Ҁ�|m��c��%�^�︰��<.V_�hΓ�ҕ���|�H����iۆ�ا���.0/x�Xm�p:aa���:�/�8b��O�O �@4�0�M#zQ��
��q}~��ǜ�8*Д�o{��L;bIF��{��HV���N>;�)D&��j�*Ym�V��,J�ňH���������방!<��	�ϫ�R�M��`��@a��ֹ�c�ݼ|=q��Ċ�z��s���H��p���,�=7�RVC��g6k��%�yn��$�k&�ٔ�!�mT�*�z��g���40	�	eW|Ç*$AI@7�U��Ch�ݤA[H�d*ITr����K��+��\�6$��+;V����
�������M2d��?H!�Rl/p��20��
yڰ+H�ޘ%6\�}�1�k|������n<6	)�O��_�FB���Py�d�*�˄�2�I�!-f�Ty��JbV^;�t�kӣ>J���?XlxV64EB    e238    20d0^ʽ�@�E���E���y W��!�
FU��W����0��j��`�������W�9{��hnI��"���(��b6����[���n�X#�EoM�k�6�po���:�Ȉ.���n6F%����x��y�=g]�EV�Y�p�9o�{	���c�\�U�äp
턮��:ԣ l�5�?�I�P��79�n/j���.i����(9�����G�K�@����%�i^f�e>�B}n(I��\��!O[��k@Y�PkE�l4�7�N���A+H��y)k.�_CV��ì��[�Ԃ�x��Q���c�r�o��!���bE��@ݽn3zE������8��w��/��㤺y輸d���Qh�#iax��,;ܮ�d~'�������X���1���e�K�@D�|I�RURSZ>�� �u9��Y
w�G�|}����D!w�������L���FY�P� zП���j�,�L�0@��|�A�Q�c]�:�t��a4�UǊ����l6�&ϯPb���P��}��,sR/�o��ğ�N�8���tE�"�!���0�i����׎|��_�Fƺ����D8�g��*�i��z#�\���g�<n'$��}��(�>HFcEj��W/L�I!�����7:�޷}Y�S�:p�@ו��g� �F�Y��_�D0b�/޲���2(�`cLq�1kF>�쨚��#�1��N�����r��7,�D4��O�~-�	{��6��$���o�6--�!�#sI��4ՙ������
{�9;�[+,��EA/�8�~4�U���9IW��.��ѧ����i5sJ�,��I��W�J��_b����B*�Z�ʞp8t�>q���6�&b���~�a�:�����~�_�����sR)��[����Rs*�-#�����}�_�[�/�ǭ}�=Qx[�/�M|R,�z�J����Y�G��i�}9;h~�U��d�����2��O@sb���^�����qJ�&*�HƳw�.�h+5�[7IC�c�	�	١p°���`����d%����?�Lū�)Q��gZ|5)��caU��AE�<fK�3YK�i}#c')(�i+~�n13�a����a7_�w�o9����>�$-��e�d~���%Z��bk�����A��N���x�[{��}s��t֡)�c�����"iF�Y�2qsNĖ��N� 2J>���'�B�(�E�*����EW^x�W�$�����]Z�ih�|�3�m���	�FF �o�^��:�)-���X���i��!�Q�M�a��wC�����w#������=,��2���K�����7���{'��P .oD�o�鉮}��{�ɇ��P[T��h[Y��T̥���VaT{߫�L��ʷ��2�f�4�ҽ�.Y�g������Y@9�����l�dH�M��S�;'f���g��� �_�`S�ܤ
�n3���;s����ү��.��E�Ww�UW3
 ��3!�'���9$��3�=~���6{��X�9�c�d��zR79U\��ۖ�-M���[�gX���P���g=�j����Xv�*�ꋹ3OHd�U`�A.y���s?�✲��ں7{O�x٘�L��3>���#y�v)�5��.�a���t�K��+��I�n2��E4ksA�'�� C=s�0��B:��o�E�����.�{��
�Ә3Q&����$�@Y��J�'f�)jm��8�h����%"�����~��������h�6&j�[[�}y�|�@ng�������e��6�9벦�#W��dw��1>��ψ��:��&��`��Y��B�6�|�����YRT��c���=5��Z�Z�+7�xS��~�."�B��d��k�f�#�Q5�J٧�~@�sE��)�W�D�Br��ߘ����KxW%����ɓ�r܆#�f�]��T��F
�x�� W��ǡ��X �j=��LQ��[O7��%~���|�0�z�eY�
lA!@�?k��� �V�Yv�_{>�x�6''�K��߇�M�Mp��F=�)���P�B�~6S� v6����G'������$D��c�\:��(R�^��^��N��ud��[N��b�I���`�qQ-�Ȣ&ՑX�����2�ÏOV��+}&DeqX��2�2T���n�m_98M�
����n�`��zg�'��k!�T���{ �Vb��o�A������7�iFw9�Ʊ1�Q�>X"#�^Z�M�e'ma���=͝����=cX����4����^D�JX�9Y2A���&���˝��� �g�p����-�XQ�3�|��z�Ih;�w_Y�D������j�ò::)�v��	�=S
�=j��Z3���`$���(M�c���wib�i"Η�̱`�� d�n�EP�/)�ц�S�Ej)���?��N��>���R��ι�pc?YK.���P.Q|:f�G
y��ܛ�nA�C�-��ŏtLI
�5�J,5�X׶�O՟��V�E+H���:��1��GxS�O��Os�B�~5�4�C�$(3�����F�#���|bd�3��er�?5�o�e؞��`�*)c��6�/a�vz�u��-j�ꟽ��x��e}]rL�f�g8`Z.X6c�\\�8�ު&?v��ڧW�pM������WX��#�Ǡ��=KS����Tΐ�>����)�@#��@;O�aXӕ̪IY�x�&���^�	bc_�Vgg���&�$൵̜�؅X�;�P�)&���\';�V$}Í�P��7C)ھ��{���,��(Vΐ�X׸�1A��o!�I��[Zz����{^E��hT2�C���/f۩��������nV�]RxH��}�����"������rI#Z. �À�����F'�g^�G�	�C�p7�q�/��č�T�K�)��S�=��.8�*�0��p�9.�N�w�M�i��nE�#
�*�e���k��k_.�]D��ON�+�E�4!�G�1�ɳ"��ў2�j#P=�I<_žo9?���!c��tb���p��7�����K:N�������Ac��ٓ�ţ��4t1�>��������F?Qm��ec�Zq�1��������ҜLz�����,�\�������Ӟ�M��`E5��Ka,���}^����8fOZ��@�=� e��⿂�^����<�&�λĈ���T	 a�hK^v�W�_���d����0{|єA%;w�r:]�2g�Y����ka@O|�o�#7�g�>�r�)}�N���oZ�2�T![��t�[PF��-)F�b�-ۖ�JcV�G=1D�b��+o��g���������=�bW�rKQ�%T�
�w�2N���O�q\R���X�m�Fx!,�?��%� +�OJ!@f�v)$�5��b���G�+�{�4wT&�%���_;v� �� ��I�)����*9���sa)Rc���nF(��E+�����l�!cx���!��$4�gC)��Nd 4.4�h��f�8�k�+�㺲�PT}�AN��P���5�:3�gU�Lͩ��g@,�zZ����/(s�
�i�)a�F�<*��5��9�h���0]����xV�7LrEle&��':�����n"�/�������4mԌ�,���`��[�GR��c�R�N+�wߚ���tqiڹtf�-r� �$�0w=�?K���ﱳLu� �\$�!�-$5uEc�>�E�8�lQ��f������w�XQ�@�IM��p^�V��t$� ��B�>,3�*����V�wh����U*��鈥��u�
�]�.�اI�h����f:pF�@߷��2�����NQ�7�0w�~<�ap���MH����̓b�L&Xnu�]h"��������	�d7�S�1.[�L��J~����UV�ϬQ=���_+��� c�b��Z�����eJG8���6���;C�[�����}�t��I��,k�h�B�g��EX/L���8���$(� �D}��|��s�In0��0�jS�!��L�4���/��h뿱���Ի���址��nE�;�_#]�>���z�HO�d 뽩�z���P��,$�%1Y��\�g% Ҭ^�_�ؐ.�f?���Dˬ���^���~T1�4B������`)�)��fL�&��vlŭ�)� ?�A�皦W�����ėK�q�1�:qaMy��')���|o��{���	�KT��t�j8��ҏ@�����M{A�U�Z���)��4�k�`dv�5�ZS�)�i��8�%��ϝr���K!��Z!L����A�,��OH�V���l�Q��e�����\h�co�x�{��M-;�Ѥ%	�0R�$߭����J������}'x���[p���`��;t�_�b#�Vã
���.W��}=qZ�M��S��Z �_['T
�n�p3hg����]q�#l�Y�����5�$�r�qt�=��b����t�\�dm���5�;��_�pN]�{�;��rg���J"�[bMo��l�O0L:p�65�^�"C
��[�fKOse����'ԉo�xr�+�>D�~<�,���6-'� �w��r��bҶ(:�j�b2<�H����Bٲ?�9��9!�m[�sRPk��^�F�$
�ذ�#:�V���/ݐA�N+˸�p�����c�졁\�N�W��B)G���N�0�G[$t\Nv�j�e��Op6org���й�2�_��W�``>puCzi0F�2�!�դ_�ź*6ݠB��\/I9\�x�;��{S�f�A�T)�luW2�_pm#����K�_u�^�Vs^/�#C�4AE��V)O[��2�͓��!����0�L�vӠ.6S���,����;µ�M�Ih�ܥ֏B��srW�3����F�(��BH��~�/�-7���d��wP@�}��B[�g�|��$�IY?4i���auGP�`Ey���F~�����Ƙ���¢N)c>udێ�2<!7׊_� �rd�s�=u@B���y�t�7[.jz�tRY�&Q3����]�����$/锪���!�0��o��|�	������c���ur����BA���F97`�C����o���ߥ��6�� W4���+2�e>f�(#�B�$x"�ށ߲�"N�$���XRj���I�'���K��HR	�P���m_�c�=jb��kt�S��B�I�tW>�-w��7�ƃ0,��S���V��)Ҁ��C��gyo1ڗ2hz5TM`����w�Wg��v��x	�ӟ�����j�"��8����<�;M��?4by�0�j��%�����B�ҖA���߆v�a�?�WR��bD$V	��)
C���bo�ha��0`�d�J/#g��)4���/m�ɞ���?x����BZJ�m]�*W��wt‑��xF�N��Ya��EI���í��0�ZS���u�[��[�w�b�0�^0��NZ��������pn��T-;f�Ӂ�},���s�p֙��rs���X�h#��&�u&�>�/ ��
�T؜�I��z��IP}SҼ���_��@�� ���4��$���r޸�@�͹9oﮩ^($�)������J@r�;���Ei������ hD�V,V�G�g� "G�fK@�$��2k+I<��Hr��M<L�~���ZL��2V���B9!/12����1+2[��9���ܰn���w�����0�L���3��� b�J�9nf�����$����6>��C w�u�����򅃰o�[D�b~�-@<?)�z+=�׽.N���G�뭜�Ҟ
�:��-<lVb��guBS����ӷqp�¼v�۸���-�o�>ٵ� �M�z���8N�T.���EQ�j�;G�����n\�	��q�8�r�1U��M���R�����A�d+���g�/�CZ5:Nc��a���꜑hݤz����$�w�̮0>��9!ـ$Bm�~ׂH���h?��ȱ�}E�}*E�#�QsD�hc$*�}�.���!������(n��Ӥ��_ɀ���,�O�l	�ecp�o"C,���٦��A�Gu
F/��kb�r:Y�T^�dn`;Jr��2�Pd��*�T�N�b��I2��Ubӕh�OP9�^A��{so��F���t�h���#i�;$�N+���'B���s��L���Gئ�id�x�_�y�"�|l�i�����;9��RۈeM�ѥjJ�*^�)|O#��Ļ�Ձ?�����O<A�:��������!��$�������}��6���F]V>�o�@����;�;R���_���[y���.����K�/��,�ju$p��#���3�?i��]v'a<�5�!��	$�Ϝ0��巚��Sڰ�UzfX�&1��J}��{�l��{"&7<�b&d�ޝ���w,�Z�sXŲsv�(@�i>�I������e7C�q�J5��D�=d�£��i~��D
��G�Ά�v�q<<	$�2�p,&�\�.OC�s&I����C+%�ϫkE��������h�?0�`��dg��c�y�.2�ݙ�YJ�� C� ��=m*k��L��|��@��bf��x��#L�%�"�V��?�"7���}v��.��.�e�fB����ٲ�{�)�dL��؎\��i��C�Z.�=�U^�ʗ�7��м�+�Z�&��u߳�
xe��?uϩZ�)��d����%�Q�ݲ��{����B������Y�q�&U���ʇS<�nX��7��f�d���ln�����'�£Tgg��.��"պ��e��[hCBy��67��/B����~�����4�tb}'[���C
���@��=��n���������m�)6u0�S�e@������3+���]�����f�j��]/˫n�����Oe���z���.Y�D���9[}mnlnբ|�͞|K7+M������p�/�����)�]�ϧU�2�z�o>,+��.�����m �oB�#<S7���U�
�E݃  �߮v��<�ac$�_�[3����m�b����/۸����vww�qh*'�B��R��[�Ð�/$9�������L*s�nmP`�����V���Ɯ6�J��t�c"z���Kw���L�ׁY�58c����Լ����	�L�Ja�;�6� {a{D	ȥ~;5M�?k�B�Μ�9Z���Y4�K��9��)�x�����$A�?���lf��j��x������&�B]Qe�Zd��n,���<��6�rn�]��z�1X9z��3�=�Ug���g̘�m��k��Z�����66F�vE�|��c�N�oz�w�D+��"������h�"����� �G�Rt��>)�q��fB�R�V���T��� H�)+����XD�:�_����/sYZ \�h�E�y�)�=��f�Z�K=2��|KEj=�����pr��S=\�t� t|4�[�%|�|�����3j�ˑ���M!�Z=�1�L�eg���O�v�JE���Nk�X���Vz_l)�����!�l<x�~
�2N��cl�b�vv�~_��5�s�l�o+��� ��3t�f���}�hhZclFNr����H�_�(=�Q�_��[�qA�Ł��}"^l��x[����di��g��4��˗����x$ۙ��h�6��3#�A���9������
�o	}�?�4���G�8�Sq���r�J�ʾv���!ZM�� �����&C6�M��:Ϳ�c�;Nx|�O�6SN�-f9v��\�����e�/y��í�}T���%�,a1a��G��/��e~�N'�/@�A(�c��;�;f��Hǁ����ضl�iA�.I���62Nw�#��a�Qi��O�v��|~�j��6Xl���p#C?A�ɣ�G�SW+ V�&�ş�@[7���=f?- ��?�iE6�1_Mi�h���X�����/�>��nDh`�s"=3",̐�M7p���M[�7�V����� (�<�;�5�iE�x��}�U2Q�D�p�} U�u�S���L7=�� ���A�_��j7��9굖�qp�����뱣�͝��tl�d4�U����1����fG�8�{��pm2���<!=nT�"�h�-�q��t1p)�ρ����?�-���"�_襰�u1�9�{���d�Y�L쁖���S�W�@��%�(d����Jx򖽦�Z��	���q=}���q�N�-���HBz���V7�,׃FO�q��@I���"ޱ��7?C��/�[,=f��@"m@�8�< �-���i�3�y+S˖F���9