XlxV64EB    1681     8a0&�jil"W�]��i�xcN�3ngHh^T]0E���4
��5��'.��&MQ�2��]���8����_P:�)E�0M#\_$D�C�r�'L�K{L�0:��T��4��lAX�sԷ-�{q�{`;NU�ӛZE���QRq<��ǽC+��#�5__)�I'+)����tv�|���S���&�#�i�Va>!�Ѥ}�)^?�$]FӮ��_@�����KD�u�0T#F��<pL�p������yVY�\�9�5Ԍ9�}
$j��E-�̄�^�,����i��d�L3[[�{�'���zPk���W�!��ՉT�U�,y�%��-@����є����Omyr�Q/RᲓeV69 �����,�"���N&���`�:���?���m��6����'�2_����f�K(�uuT'_<��J����O�r�z-v/�%�T��1�椥#�*Ǒ���Ͳ@���Y�V�DA]\�\n<�Y��S��H�!S�Uذ�

�j�f`��KO����j�Y�a��؂�O�bֽ<��+����,��7��븜�^�Q��Y�������%��}�%^`oa]l�h4� E���?J6_�eͰ)/T��>,���s��ejF!�D�r4idS��W��ˍ������|Uӂ!�t�Y��{C��Y��qK�����B�OI���~�2Sz�XMQ�,w�1jBk�ֺ��M�o�"�.s@~����2J��f��mGf�҂�؝F��N!|��p���p��2�A��Bq��"2<�P�ۜ:	e����G�Ӷg]M	�fOnG��ZFS;O�R��ϵ�9��t(8U�+Y��͜� �%����W�|���O��#�pA#���;4�c�q��#���(-A�涇[���h��/�p&�f�&�W>���/l�1��Kc{�	5�'4nW԰�y��ğj�>4��`��ґ��N�՗����ױaJ6 ��d*��@���'���W���L�f"l�K�������@��[��r�/+���w����t�����r0��Xjrgf�M��"|,&Q�V���x�ӿ,iy���N���eT/֑F����wn����0Q�����.�Pͣ�T֋�tq���	t9��%�ͣG�G*���"��8�T�g�	rm��B-F�e8ft�n��B�J�W��J�/�K�2�R��jV�����K@�QS��0�W�\! �������:ٺ��A�9s���t�+@��*>C�1���މ���44c��>۱�d���������D}t�bi
y��%��W�w�{C������p\��q��~�#�!�m}�	��,���Y>�re>_Bn�𥾰Z����	��k�����I�R����P(F���,Sf;gM@<7ڦ�y��0�B��ݨĐ�y��S]h-��1���W������?�|䘽 ���]��~Q�^����3؃�ȕub�͕2�+s���;a}$�]~T�B����m�Z�0E��sm�;i� *��*�H�s{ ��;�#���]���4���Pn�"%m�H[b����3�1��+��:g0���*bab��%"t9�x�������?@-��*f�7���.C;!+u�^����W��p\&��
e��ұ��H3G��Tʠ(��+�8?B����]�6Hz�m_=x�Jy��+��63�4$P�@7 �VP�ڃ>�4Z��[܎�-є�21�0$�^�4'�^lC)���k�`����\F���Nq��ܨ8iPc����~�CK�aI�陯i�?�\k�#�C���4i�w8����9��[w��������L�D���2P����;�4+�G{4'sVu�C�ҍ��'Y�&�[^ê����P�i�D6�)��0j��)sU#;� nvC�\!���rICꡔ�	��W�F��|'HW�������8��愆�:�F��{~`�
�m�7���1�o�9B��ǭ�yp=�� �
����xB�p��H4L���s�0�5i��k} pcx�^����>�<��!~����O&oY�V� �6J�J sۇ��%!�A�B�-Pd���L"��HL����f��q[�%u����k���1��;� �SF�ZY��b!I�JD򇝅�S�Md��-��(�YȜރ��
��`"'1����D�C�E>��I��M��