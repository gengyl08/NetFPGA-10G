XlxV64EB    171d     860������g�7(�{�+c�*��wc������Ki5���?�17<�_/q�3.�XHrj�@�/�3'���*�(���{�p'x<͙��{ڄo�ͳJ�G?mYw�c�)w�L<�����c����;��m��1�,���p�S#�"��;a���"�mqн+!�ü���U[�̰�?q�L�Y9�p�;���������h1.E��!rʖ�@�H��n�1邤ň��1�"eS�a���N�e���1'Kb�r�� VD�lZ�,��X��G;GSc��X���'��a�M6%GX`�Ͷp��La[I?���0��-Ӂ]w�	�����KӃ)?����<�X�̉����Bx\�j��H=���#gT)#���� I~B�ٺB�w�e�͎���.�ƍ����_ �^ - ��HK�FsvV����.SY.b�v�+>a�|��PaJ���pn��;��6C���,HF��-�-̌��T�B�A;�:���!�Fu+ߍ�������k���R�#���w���_v&���1�(��!���<�6[m���^���RA|���閺�����N�e<uq��ơ����8؀�Շ��}�@�?0���
>��p�~U>��z#����u���5Ź����E�UU�fXX�m�\�����m�����
<�]�б��,!��~�	a��>4���ۮ=7���?�b��{VR���	NIx��h�D �g	�y�6��,q�r�|@;1�ެTWFNKd�%���J�����d@6���'�i&�������/��
���`��>�c�aѩ-��x>X��(~�b`S�$�C4z��i�e�L�ulUe�5�X1k%\"��W�x^-8��Z��Z\�Ԕ0F!�2%�:dpl=0�&F�?�h%�`K��EAJ;�\$5�}uZ�$��c:Q;����P|>�4OeR��"���{yK�D]�6=�^�)�3*��/�:��$�9W�j�Ɨ)�H(�xj��[�M���YdEۯ6kACԃ����v^i�� �F�eS����eVB�'�۠Ã�*W?)�����B�j�w8;]2rRh��K�6��%cG���J`Ґf)��d���'0M&^Dox@�fe�y�>��?�΃�{�x�o'�EI��nP@3��؀�?g�F���B������Z�%~�t�Ғ4)�iI��9A�����B�D�4�*#�j{IWc8B��F-i8K�SK��y�%(� ��{�	�{�k�!�8����:��2>з�c�ɕM�p�ʅ��}�7��)�/!#Q��mԫ�س�v�t���t2�F�#��{�׃�gA%]��г��`�,��7�R.�}_:!e�v?[�S�-�9�e�v&���])��,�\���lA�J�4�a�]r%;��J�/�]�Ӄݘ�����1H�H��Q�,|$��`+��d͇@�E��H�a����	�	�b�~j�����r����HP�Bق�s����];jATE6k1s����Y�K$T�:"<$�Ү�z}��U�t�.���۶�&�>��7�3|���PJN6=3���Z���S 0��H:7XVW� mZ�ot���i������	"�J���U�c,���EZ!����P!ۯNd,�ya���(0��� P+���W)�"���߁"�pt���vn���' �b`���3%�;e;�(@�.JRoގ�lc�G�*O��r��|����G�����C�?�����ŧ�Q�	�(�����m���6�A�.7���h������4}��cF�J�)i�t���M�~��8@\H������l��Dz��G�q�t{<��2�I�c���l��=���Zr�
Q1�6�3-h����/�Q�� �GXY$�4͒y��i��\{��|���{6�m`� Hh��T3�\gW;!4�9�����HB؜�B�i��*� ����'�R � ����>���3�㓱���?�7"���J���m;&���+�$mS���藫�u�������U1���5(�fIL�t7L���t[�y�I	3n¡B�.�<]��W,�n�O��֯�ԸA���o�MK����De�lb��ԓD��zx5��C#��