XlxV64EB    2121     ac0�� JS��࿫k<��o�Vq�c���,>s|����ZpG��s*6J��x�����*}!��Sz}+y!*�0aa��Z#/L!0XKĪ��@f���7�� ���J�X��2��
���ѫn���%���G$>�h�����u 6x���ٶ`�)�f�E��ͼbn+��g:�[��_~m&��w��~���;+*" Q�<�
35*���G�s�?��iQ�e��c�-����2�6�,\zSd������p��xT�q�]�?(��[\p�{�J�/
!/
o-����gX\N�AU��\�Z,�I������H��(��ziN�{#�z��<�rtL�	�Հ��Ǧ!��,��ĉ{���햷�	��PJE�{���ݣ,���3��� X�S���E����E�f7�Qy�(>%b4�}5{��[��)���

��AU����c�>
�mHFkx�X���P>)��c���;��
*z-��tjB9�7�@s��lLnx�j�ey��f���_71�#�ё��m��:�?�Q�2�y���rfoBo�+��M
^\A��M��Z�70ϼ��[��0oq�+S�~���1������<�{:�
B4=eK����Kj����+�s��?J�5v�1�ԣ�Ur�b��ӁN�uYqE`����{1��5)����\<X�qT嗈^�K:rd�Lm���j���5(�iA�r���Er��ͽ��
Jb~�!�o!�k�o���	42p`&�dӛ�OH�VϞ�����O�v�N�4y���f�]��d����7��K��)�B�	*�]:�a��H��`ն�gg�^�� 5�Ƚv�V���ަS�bZB"ɩ���'�Ϥrr�W�l�.�I�[j�|����X�Q�%�=3�z��p���3�BL�p�-����g�XC?,iY������
�+T���Xw7xp�oƧf}0�-����Ü�}����ٴ�C9ǥӡ缃�"(̆׶۶���lm���\��U�
�>#�'�0�B�V��.�9�9`	}-�>F����ԭ%;����J�vu��"�ƙh"�s0���-hVuU�
o��m�W@�C33gѠp w_N�5�� �K�g
���M�f�5�Q~ߨ�ĔU�nH�e��0�l�v�ƌ�T�M�]AJ)up�X�̥��Z�\�@�#G#ӄ��[̤�䉮�bC�e�;�_c�U���"��U5t�'ȳ�\�W�?(H� �
;3ͩH�2�����D%��\R���]��	�� �<'���y��$x�Rr�qT�A˛}�>��刍� ��E�&��sDd�{k����1ߌ�ڢ��B޲l�V�h�-c�%�`3�M�g-}��e����P���_y��	�f}.�����_A�,�PB#Mam�/g������3Q|��?�>צQ��ܤ�g;��q�ޞσgc�����0qc��L�)�뽩�(H�#�4�*,"��a�)<kq{D��ˏ���-k�(�?�}�O��i��V�f���j,�z��?*07�G�!�$=��k~C�%��[YsԂm!��2�F� �����)L��������Ad��A�o#iC8Ir�:�"�-w�QLV���������u�8f֙��֥�G�ײ|�����ٸ	+�2RJk�����_R;Vw�ܡ��;ÏG7ϛZ�N �K���Vho
_�5��=�.�;��M���,tT��!@+���v��<�b��=��',�#%�B�$�nf��b�_�ʐD�[��z�)/(�ݧ ��/��)C�������Ot�߭�I�<� �EA?�ÄŨb�&�b5Q�;a���.�|��Ś�7�=�ȡVu��lE�'L��+z��W����n�)�n�����!b�� �~o�E�{�cר�������I�QM�:�������q�X������rY��P�_G��y����R�4r~rЗ�ı�0e�T9_�`!4���&J`��N�+YM9�Jӑ"u��ۍ�*܁���^��l�Y{3���MK�-�,���B3:I01���e�� |����7ɕ�.|�Z�[��˫a��O�,U p`����K�@WY�J�A	�te��4�P������������_˜zɾ�a��>��e\�O�P�|.d�Zm�=3�2�n�~͚'֪q�v��<J�e8c(��z"=^�VA����(�{9Lf�[fb>v��3���r��Ŷ_-98��S�W��ꗬ������홠���N��]��n����p��>^Ic	%�5��k]ƄN��z)�"�o�_��6�Sf�$b����].8�-n�P�I:l�;�ȓ���<��d�Hm����oV���.�w@�-�s������҆�۽��l�d���ع���A"�D�Ռ��E��I�	�e��%�?.S�7����;�E��Q�5(�����d[ֶ@{�x4��_�sju��*M���N$�O ]V�Ҫ��D�!�6>�ޑ{*�`hHSb�=3�r�Ka�|c���R��1W�d  E�C�y��	�.3K���߹���}�wv1�W�S�m�b��UU�����D��kCLd��F�	�O���``���b[����q��0;��f�P�'� I`�'�H�-*��G�s��n����,\�p����~.}��������J�K�[Oϔ��"Z�.i֗ �7��d�<Z�؞�Z@-yg���W]�+w��?�����%��"�?�*�bIʫ?}��