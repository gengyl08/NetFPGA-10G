XlxV64EB    3eee     eb0`������;ti�/�AB�b��]�c#p����fk6�r�~U�B��A�"�H�5d,������l�M����4�]'	�|�o^D��d@����v0�aҟ,"�H|��a1��Ɍ���v�{�X@On��M\���87��C�v�v����d{$�����"�Ҕwzf���c1X��PND��?�V���,�Վ�㍲8��� |�B۰J�N$"�>01כF��ӑNCAҥ�C��_B�x�DR�K�u{Ɠ����� 
`ae@h��$� !(��3f(�xDv�7W� ۮr�tQ����=�V������1xbH%�`���Or0���3/识?�U�Zº�R�S�\P�g�7������pv���8A	�̾SM�IEs)��� �gF����XK�ᴅ{����e.��X(v��̮�5��а����/��� Ȁq��K�n�|��R��N&�}�^�����p���"�	��|�-
#5��b$/H�CR�4N.�h�TWU�����U�����p����}��ѷ�NP��i�gNy�ӑ{KbE�8�?[+Rr�?#FA����1PGx������B{Bq������F9���ݕ�@�Q;?����i�s���	v6C#R@M8EJR&~����k�Q< ��?4BJ��x�9�y��f��EL�M|�cim�T��囧i��P\%�Q�]�m1���,�;�>����Lk��}V�}����c}�,l�(5��F�h*vH*<��S|��7��$��l�@���ħOOl���;��P�!3��J����53��V~��]�Z��]Ȧ&�Cc�U����٦��Ev��u��0�2��,V�w� F�����Ä~l� ;r��r��cӄ� ��ټ߂�-��)e�|��K�zC����=�� �9K���r�v<�C�&;}���cS����@�L>�O@PX���=�b�]�'��y���)�'Cl/��&鉤�]����ؤ�݈�%(��s`<s���PT͋k�&�1�cG"�U�᫪�?MγχSh�|*uW�s�y�4=��@7��	}ԮR�1ܔ�ﲹL}�Ĭ��#�-���"�.E{>=#3�]���h �^�]�Q�);�.EC� ,	Z����+�P�r������n�^o����!`;�.u����=%�VҮ<�c�]X3�q\�X~��?����+�}���˩r�P�ݩ:�$�^_��� h�"VV��ݷ<ǵ�S�+�2�b-�*��r�~��ܴ�Ex
g��=޳���o�_�7���W�If6����� &�Z��Q���Cw��Q���%5d�ख#86�����O�H�xU�V�A�p�b��keX\��MɈ��S(�?7m{_.�;�O<������|%ǔ��o�(7�I[f	X�I��.�(Ycb$&�b��N�˟4��F��Y��(�1Yd��K��2hM����8	\_�C����[Փ��B���$v'�=/��������v�X�G�>���̂F�`��4�3f��j�'�����Z�5�?�L�Μ�%����r4*>���[M�&�'��&��7�#����%��Vr� �Y�.˹�ϰ��� �O�H��?ג�(�eg[{��f1����jH$����	�����\ݖ���
X�!�Δ�;4�t5�l�iP�i0�S��VVxSq��KQ�$���T'Q�'�qA�gQ�f�¬��o� |��V��U}A�.�\�
�h�+����q0�V@ñUd�� }MY���u7�C��ӏ��a��%,���Ä�k��uo����pJ%�S��w��c{w�b�x/:i~�N�g>��?�K���S�^��(o<�Y�1��#��j�R��H�O�Peش�gR�ȭ���@풅e�s?�~6�ۖ�^5�I[�}��`� ˂�T����
M��`��<��� "�Y�)Sym]\��
���{<�������I2��*���&���$t�WmT�t:s�7�owT��V-U�]법n=]�1���e鴹�zo�M�X{қ��ۨGvЃ���#����'-5��.�h�";�j��a�<�J`b�0�<!{�|�W_(gv�#
�Ռ�=��3��`����`�ᐈ��<Cn.�S�����A2�t�l'��M7=ZdҠ�����m:.���@3�߮��L���=��k�VC@g�/�q�p��*���x+��`�1�=�~����O�{Z��1F��d'�f�=P��BY8�o��W��'��hk/�w�D	A�*�L-�&`NeH�{�x��fJK7ᐺ�3d��E��q�KI��)��@fH�"��uo���j	�ˆ��
�	�fE��H�GIn ��l�-8{B�!5�H��Lk%�֔�|�8�8��#��4�@mf12z����z���Pd����{��	!O�M�'��VڋT�k(��v�~��C`��7��h��.�F�Y��Vב�'Z���55?����ʧ��h��ɾ���������*�K�J�nX�\� |�s�3Cj�P, �%�p7�[Ġ%��xw,Nmj�^�F�@�=�{l�����z��R��"S~���l�'�T��ws��1�,����e��%0� 2�_�s�O��%�օ�%��2f�[���dh���ٗ鑌�����k����`ȫP���+�6�!t^v:��=X�C�ј���j}A󇟼�O����q���ȇǍQo�<JA�B�;p�2.���fe�d�Op]hfUT�-DC�t�����W��(�L�����ż����m��������nC��9��0''���{܄BO\��"Z�o����p���	���2�*��ps�gQ٫�#gw'�GQ�ur��\NwM���ܿ9P�3���ć�յ8��p?����juR���7������65J�q�ݙN�9���LCE�&vŤ�?eJ}
�z��Z-�Wv�<���#��"����T� �-I.C" X���@�<Ϸ��_P��-�_aɞx��g�V<�m©R���_ad!n�Ɵo��6��a�8��N��B�h�� �j��^8����zT)���U���G��Ђ�w	Ct�g�v�m �&��2�[6 8��pH�so��ֶ/�;N�O+1��-��4�t55�,*���N2���˧�tsܥK%��ľ;�	~������dS�J��:9�� JB�B�׾f�����|r��=}�;��+�_l�4(�����nyצ-�|��z���g
���)��z(Th�7�G�&vCKo=�����5B@�˃1�bz�2k>��6#˛I�G�v�����c�-z��V]��ȫ�1'Nԁ9��A�<���r�*q���%����L�C���T*{O�d�:lK%�e��OBR�L2��Zs�����sS�Q�nw �ؽ�=1~�a����_������A�*��Mx�v�m+�ql�
���e�&TK���"��f�."Y�g������ g����t���.�&�el,6]r
"�ZJ�nl���K�s���1C^��*�h�6B�{��-��)M Iy�K�~�?����셅���"l!�C�� ����/u�3.u�,8�6S���w���g)��Ń�F���r�Ɉ��F�\]�ɹg��|������M�	!4lX.ʥ[򦆋�������`�_L�Ii�[�@�Ԟ�"���Ƨ�H��A��}���9�Y�-�ht�e�o�*@��R-��T8��K��E:�