XlxV64EB    fa00    2fb03����x���h2�e1w�cn)�����+��*���v.��׵��ε��P3~�7�}�+�4�m+{�L��ٱrdc��K��d
�������\(�����A�Œ��ҊY���Ӄ�]��&e>j�dL���	G���\C�Vgs���A�˯.&��Pdݓ�]�d֬��ĵ���h�S����~� `{ף���f�R}'b�;�"�މڝ�E�gf�ӈ�hR��=�X�<�8��K.���5ڸ�5p�3&�)1��1o��G&��C:V��!�?�"<��#_Gs+5�i�AxL�9��ϽUN�7ဇ��/�_��3��������ة���&��\�[������������s�d��xSZ�L�u�4`<�|���]���Ђ�zu��"f��:�a9�ɋ]�\Y4BAy�TDk���x޼��r:����+j��d����&��cX���9��z�8��e��
m�8����������'*0e^d
���˞�������wxtS��c�r� � ��k��\��m#ّ��Y'��t7K'p	�3!f&����k(� �T�x^;-��@;�D���=��k������0��Q�r�s��m�h؄[g|�����ݸ��G��Q��@��>&�kn�B���,�T~��tӬ���yI���êE&�L�>���/a̸����x��<�(�Ǵ�n��JT߷�Y�������~J�ٞ���7�8�K�TN�a+��l��M.�߶ػRǦ���*v� "��L@y��b�y ����ű��AY�HO[�?38+K�Y����;cL�I��A䪞q�~)Ki-iO���N��J��s����'�|\0� �ϛ��0A�c��e!�	4(1���w�c��4��	��ą�g�Wc�q�?�s]{�o��q��Ձ7ьM�w@Q�	�<�@6����35U�>=�����tF2�Cɗ�j\�miO�\8o��E�����i�p�bA&���^n&K�1���N��f��M��J�@�4$J����x�����s d�����$����e��'��8 �����g�H��+�T��Lb\�.��z��8�/����I��5��W�(���� X����6����^<�B�)u9� �fح�@�E���f�g��˞y��*[cڌ��!�*8u��j�ؤY��Ҍd-�����Q��-�`�YOS�kp}��/���*�4K\�*qb�jѓ�{S�<�]�"�+o
��[ w��d�lU v�vM�	�!�0_��2�ے��?FV뿢K��r�:H���_t�E����b�y:��jF�D�<��@�9rƣڿT�#��H��w�����RЗ��#�S���a�&�b�R���3s��#��b�u٘�J�EG�A����㥑�h�ж9H���h\:�xefJĈ�.Pϲ^�x�Ghޔ��́��j� '�ۧn��tܺ�?�+���Q��������+g��!\ЛK�L飴���v5�05�H���(����c�uU��U/T���}ق�q����ĺӛDP��r}�_��^]<.+iR/���&��E�����C���#A����N��0M�7J佪o��}�g@#2�-GF��ƣ�ճ)0��\���� (4�:�1	�[�� ���U�W�=rWH�AϵT"�U}���a���D<�unmZ������{M*�c3�e����/��;�l�/�?�`�Xbr��m[��vozo/8��O�����ŧ��C�D�ry�RY�F���~��{>u�ó����8 ��IB���0��^R�ɇ����5�x����hc(�B�D�QQ�K������"���(�o�����I-JF�ʐ�n�(沇h/LS�����Y��*�~�1�5��m�����G.y9�Y�>%=w�H�㦪5=�R�p���Rj�p7��4k���QAR�8��ב��-�:'<kfq�����m%$ER��Nn��'��^0��l���r�X�Bg�e�z�Y��Oʛ~���b؁1|���GY���}1E\��\Y>ɡ���S�ŕ���Qa�� >�.#]�g���U���(� ��@<�s�e~�}n����LQ*U8fBI<t���p2�i��w)Q��&�)q)��F>ɐ��8>?�7����l	�&��4bƶ��X�xh0��ǿ�u#�Ž��D��%��"+��:�cmvl;�G$�
�������O�6l:O=����B5��}���e��4쩦g�
Ѹ���^��k�������N*7a)ޖW�$S�8�929��R�GgCkٵ�Xև�ʚ����弻��cM�i
�X�HR��}؛�^��p�C %Dl_i4�n�s/��>V���G�Y�ֿ\ZR� �c�s�QP��I��K�E/�H)t쎠���ݶ$Yf:�Rt���X�^2�l�7���d�"@u���噾+1f%_�D�
Ǌ�Bw�V�'�t�@�� �!�u��Q�Bx��|��oY36H� �������z\"�q�B�/i囩7�}Um���f�vG��>Q�΃��&�16�*�qb�C3Ǔ��8�^�\�`h��|R����ǟ��t�ݫ�����RXO)F��_%UJ�B�M�F�"2PY�B�'�k/��a���D�'L@��rE�����ol�_��"C���4�@Za�<���[����R��=�|n�}��?���es��u���Ƴ�fٵ"Y-��f(̴P����t]:Z7C���A<ϋ6ȳlGa�2�S�I6RI'.%ugj 5���)���0�����s��(>5�BgP.�Oc�:����l3����琇њ�N�ݳt4���]3��M�=��t�������"�����7�:�N�&�'���S�llE�k/p��U�/I�%U~L��X��ߝ�k�tJ�!�r�����`�?��~�RUT�����;�M�0FO�ť:�~���Rt���([�NB���5�n)�̩i@��%kE��4�$���3#�q�VYH4������`��rx
����U�Ġ�G��Gh�+uK�QM}��pH�����Dt��@��w�3���!�[��}РHc�}mB��W"΢&2wZX�#c��\�p�����T��2	[8!�rz��Q["�$��V��I����܃��R��+2�R`Ҫn;����z��޿pJ�ރ�DDO��|�Ԃ��_�l��z����f��B��Op��J����=�^��fv9��~ryXW":�dDBV�np9d�����p��I|����ߐ��8�6��`d�K�&,���O/�X��n�Z	掶RRW�0�S�Y$֠aω	�D��t�y�,�������iF��;�gz�Gq!��Ks����ChTD�K�/��)i����_�3���	��A�/<�V�4nS����V�P�c�͸�0L���Yx�ܫ�ޥ]$��\�]Fv8١��ىn��7����eXn@��Lٳ6�\�l���kд�l7[2K���]�j��x������
�"K�Me-C`�� �����F�k�H��t�v$IWn�?i�
�BǦ����r��[�5[�_��ϳ��;(�/��uo%)�sD�%Ej�'�0&��a�T8�����>��2�gq���-�tIq��"�8v-[�Қ���a�i����\��yج�nbx���O	1I�p��PH�H<Bɜ|m���Cu��0-N2;>��B"*�����%�O:e�8B,���s�?"le�;��/5;RZ�ƨ�K�׿dkS��]��S��P�(�+!ʳ��[t�D0Z��iΌ)�z�^t@4��(�k1����9��H,����� �Ù9��jPB��u�P 6�8��_�E4�1�='_��2c|pa�TUkH{G���[H�ò�Z��e�2�ݑT�4h�`~�I�ί�E�︵��Il�;t�� �-�֥�L�����,}����x;�4�1�n!�Ƃ���'p.z��j�^��^���[g���gԷL��x��-K���n��q7C-��v��rQ���{�٩k��E�v:��B�Y�@�MoaoRrp8qX�<�$_y X'T.���{��#R�Hizk&��`bMM ������g�Y�.�N��w����
�c!^��zC�A!�� R���ԅ��!	\�K� G>�=��f��'*��B�V���;m��O��i�JzK'l=K�yO*ck�Q��
Ҕr�x7�j�����|�t)^��ԝ���}�H`�d��+�����5�E���c���Ļ~�|�R�K�>����! �P�X�rv�9y���x�ɵ#��U�P5~yƥ���7Ӟ]�?�����5�*t��M?�����!��U7:�(�W2�K�w��i�'*�[�Sù�U>�|.ۧ9x;u�8o銆vQ��q�Ԗ�[ep�!8��2>�"9�Ks�l�͡�Т���?�5%����Ҁ��u��K��ګ^c;��ip5*��`���dG�{A���6�&���P?�^���r�Y�szZBѢ\M#6.� �7��ӛA�4���X�(����O���u�w�F1�B�A����׾$|���X�gr��f��S~��|/��{$�q���{���(1���&^�5����זZ^!�KxV��@y�NU,�TB����s�>AV<�Y+ �h��QD��4ZIr�s���Ya�!��?t~D=�,�Oǅ���E2��j*O\JZԭb�Ϻ3'ǹ
z$�$b�Y��x��;���DNB�5>��Y3��`�i,��
n�]D/��_���v��ƵY�(i��pk�GGD�n��rz�K���t6�RA���(���6��9Z��%6<�8�p%Y�������;_�J[�Ide�j�A"�f�����o}�{�c`�	[�&c3�^���>���U��$�(�7��9�\>�Ҙ��~1���:�9#L��3(y��3x&��3�4���n;%�ĮS�:~ })c�~�џ�G"��+�p6:7h/��	���4<�:I�i��(R��<�lU�ؚ" �,K餛��x�S�AӋ	�b]�y�.�Uҭ�A���ܭ�"�ǭlL]�HD#���Q0�]
�Br��kk�e�:�Pn�n7�>�������C5k@/p�d,����m��O�4���h��i��m�G(�<�>��v2��8�{u�ʿ�u,����j%���LaC\�i���Y��~�8���_��S
I��K����ܮ��A�v�<��һ�����F�o�4�"Vs���ؚ�P�.�A���eν�CS�>�f�U�LD�=�<�t{�L*$Q��"Lj~�Y���i����=���~��0�y��[�ش��v�j
1�I�~n�(���M���I+{�%|c(*j�<[
+7Y���"d~�,����-�ޮ�p�;c�-��_�ؾ�O9GN[�Z�e��Ko�58�G��'_�dg<�%��߳�4�����ug�BHz����$K6���� D�r�� j�x�~{Q:��67Q^t <��ve�>����O���#��N��a	+̌�9
/�!n��I������/�g4��y
�;�2Ҋ֜�{'&�/}2� ��p�s��I�{��(��ܢ�;���La����[�,�Զ�$*h��Y�x�C��j��:��ٜ���U�=���Lbx��=���1��S;7��?��U����H�zf��񦭡�������cy
=H�A��UA��l����ڕ�i��؀d0�h|�4f��r�${4������!D��#̣����]������	-Xꌂf�*�?��
r��&���+�K�=I43�F��BA�޶#&�ڬ���9�Ƨ�Lt�zG?/��u G��}�C�S�g�K�icq��Nw1Y���F�	}��i'V�8�Dg�礛KT�W{�܅���"�)���h�����u�'�Ԛǅ��+FJɛ��Κ�c���ڝ�R˛Ax���~��5���O��NÓs���b7��2	i�W�D�e�-��%���%i������͓~;�E���3 q/�?���"u��)�D��L��6	��J�q�u��#TV�Ɍ=�GJQ�Ey5��@�MN�����]��g-|1:}V��e�h������_�@��:�P{�� +�J�: ;v�.��qx͇�iD��!*�. �b,�B
�!ۥ	���+|Q�[�wP�6Da��il�z�{I�p��ˌ�瀰�=is��7ֿ?2��^�L㏇��,Du<�W�`�LZ��h�=�_a�bj  �lc�V.�|�(�Zm9��Mbr�����3j�9����$�}24AG�F��V��
�H( =���
����6Dq^�Z�}�\;ӧ�/*�~{��2�$�B��1Īr/��~�.}l��`�y��4x&�_U��a�1c�V[19N���X�������)c*�Ȑ<�@�d��8%D��/����A�wϙ�����	t�ʡ�[�5vя�z���8*����bc(�U:�_�0��,���^��Xݓ>�Ԕ�
?es�מsr	!MiLӦ|c)�s��:t6�	7ZҚ�8L�RQ������ʮ6�*��P��N?�Zt�A_�,�E}��W�!��e����14��6h�ss��\=�����F0|�8��kS.��Hfu�{nnY���3�Y�f{�4T'�)B�m3��R���[X%�B�T�o�(�X�.���>�_s�43g����ŨX\����<]@�$X%wK~E�3�������p�_��M�1'!U�S˄�eu�;������_lf�e.��[�ž:[g�'��6]갋L�Ě�y9���*�#�;��bT?�*6�Ehx��oΚ�TP��J���������C�,��[�$V�)C��N��i�0 ������V���dQ}7��gˑ-b�-���n�v��S�(���+1հ�dBZd�����FY�mROl�4��	]�CZs>h'���280w�SIR.�%�*��sR(Q��mZ37�H�z��d��}�"t��gk �e����� �r~=�+Q~c�x���� 0k�tQ�\K���P�����hB�������E;{w4	P�J��US �@�?�򱼏Q��t?��?�����P����o��E:C�\�Cw�` v�V5gz�5x�k�8Ağ��vx��
�J-�� ���T�U�]-�A}��Ǥ�x�׻Y.A4	�Rb��1��O�b��P�ў�5YB�p[��R����]����6�CH�d�QCy�N���]��M�$��R���+n�F��mɢ�Pݙ��	\P����B�g^��]�R.�`w�y�o�xw�_`��+ߺ�Z��f��i������g���S�fijTs{�
ۓ�!aq�.ni�]��\��(��8���"�����-Aa�R8��sy�s@KƄ$+ESo糣]Ra�fơ}H�i��=$E���o1-���j�0"�Ĺ����Fx!�.K�
�C>JaĲY�Y)J���Mp�e��� c�"l�m���#p���+�t�2c�T 4g��D��չ6���}�$�/�Ap*ilwdǾ�5K���#������>=�9�����;.�����6�ͺ��v*�Ȧ�_;M-y���SW�6_tg�w�]_��)Tƾ��z
�T�#��zj��,Mӈ�@4����Ʃ���~Jh�,���G�Dq�h�`��a�(Oΰ�h��v(Ofԑ����8zܓ��C���[�Y�V�w'~��(�g�A۩�%�Z�� G����<�K(v�qg("�������HBH��㙓�p?�7���Z�� ���u)��+)JB�r���m۟�*DB�[v?4� ����=��ri�z��k�%�s:���+c�y�%A�5cHiϠSl�wM�B�#*6��Y��<��T��}�-��̀�����ph���"z�Z]B;�v�
��0?SF��5ؠ���:�����<�r��v��!siE���\A>z�cR���ɑ�)�Q �9@�4���{,�$�n��"�x�ޥȫ�2|�~�FvLl�ud��N���c OkSK�i�
���.V��:��c,܏�P@{�F#?2���+X��rc�+�8�V���#��g۲�o1��F��
�6���,Z.�=y�A5��c����G{J�)��WT �:�F���B�La�̑��z�BC5;�A!D���Hr�E���Ȳh���u���I����ܿ���߼��)L]�F�Qo���U�u�(���z�d�RL��;̤�B�,�2��H�s�f��q�sK�[R�~�@[}gٚ�-��n�L�è��F��4}=CD����;�o�����;����DOӗ�ץ�ۘ��1�pH����˲�}����	\���������d�zr���#-�$��%�T��ѷVW���F�O�����@ۜ�b�������54����Rw�jP|w1>n队c�4b�vp8(�gFH��[�$���v�=�1g����07�Y^�����	Q�5f<��Ex=���V�I�Ͷ̗�5�˴Jl�$M���:�W�+9���l�~m&,
��7��葕���[��'��sTR�N(ЛۯH��*�D�@{w�!��̚?\����4�5[eQnb<����+l����o̒KvB�"��Z�T�n��?�M0��-n�/����il^z��ә��xZ/	�R�������l���*�K^'�;�,7n�A����m��{F�urٵ;��M����5z�" ���5C������W��N(4�=|& �0�*�n3?sл��s0��{��q����QYR�nʊ娷n�$.=u�"��&��QT7����lwg�a�E�P ��y����̌r���_9��U��uz(ت��^�|���V
	�t\�+�|$�YQN' �b�8#��27��u�����������3���Y�?�}�
S>�|��5Q;p��@���k|�����.��p��a]��M�.i�es�UE�eP(���f�,�uc����XEA�b,-�2K��G�����P�J���X��y-K)�{�#���r�X ��TX�K����I*iXUq���Ut&���0��K�%��'���e���&QH�������*Uf*6���{��G�hNE�ǨM?/�C�kyM������v�������-�$gy�a#�����7ǡ�{��Q���Ƙ҄��1p���"�q`�i�>���ɸױf�WrgIx.���0�^�,��b��,҅�v�[0Rz%T��
,�qW�x?���
����*"-N��B{�	�RF����-"Ζʝ�&��g��0~���2A�6�!ƽ�)��ɤ��� ��x��2��a����\D�τ�͸����ꯆ�\��{~������+�e���ޒC�)�-3���ܣ��!��R��58Jj$�g"8kA@o-����_K�}�hX����K2c�U��-���=�;_x0�؁�و��޷�3(��[����b��Z�hi�_[���N �
(�P	����},_cʞ�hCy�џ�����òj�.�f��/z:� j�5�wI�e����\�\�j)ϰ6��W:=��:�-�^���VN�BR<��e){dZ�m������m�>�Z�3�u��c�_H"�����@�T��q���"���aB8�6勤��W���/�f%�6f�zH^��.��]�$�3�?����?�82�@���Y4��]�ߢء���#>�_/��d�����[�;�T*3ܿc���r�`�ֲd\7ޤ2d�6��%������@�����y�A�,\�fb�����{���(o��]J��5�Ǧ�$�����p)h%���t١+�@�z�*T?H�1���3 ���[� &?`^�0�����k�G��C�S�	��Լyr5=�q�HC�<$�'E���سCM^�b�+��?��
-����	4�(O�z�������_������7��/�a��|�'����A�-n�S�-�b�c��v��m�k��\��b�А�j@%�opkPW����5��UVЃ���]��HhC-�s�;&�[ҤPg����Gד�O�N2�y�m}�٨{�4tnT05�5$�G.�JF�s�-2��@U?���I����!+;�(��-�I��mv��Y�]`��|�a1��o�6� ���?و�J�+��3�7������+�l�e9U'��0��Wp�Hu"]����d���X#I��/kU�)�U�m���3�l⚗�1:�*�lN^�S����s�5��_ȑN��C47Vw�z��c2�����L���Fu��V)�y��+�lt��#04��T�V�k6��;�0'�i��0�P ڒl͚%��d��F��YZ�;k��s�F��k��ڹZ���
�ؖ�;��6��	Di�x6-����i�k�M�[�/�;{5�H.-۰��h�I�І�� �Ӄ��/�wa:����X�aΒ�15pK��U[�rZ��W"�Y2���'�߽g�kF��"a��}HřM� ��I�g�!
OI��P̹B��ٴ޺"^PV�!�H�I�e��gV-�u�0�6$�aխ��M3���O����n�A�_�Z����<���c�Ҹ�[��38��t�H@�e�%�i��b���R�CF+���֙*���YfIl�r>zdj�֭򲝾�(t�2���E<>���I�o���^i�R��$��9�������0�¯���J�q����c����=����P��'�W�£RM7_mޯ]@;�+w�Ds�ZVU|1�?�Nq^
iO�f���̳mVb�^|��1Q���&āZ�-R�ș�_�#ɡ!���#_,���N0y>ȭ�˞�p ��{,^V�jF(�4�����X�:b�#�$:���IA�|��è��r9�_B��|3�"���z~w �c�`��T��B�4����)ȍ�1`Lf�`jDSq8u޶b��o��n����?�/�<���
�u4fЬ8 ���0u��E��)a�ǆMn&����m�
�3������s��?<8��g/@A�@c�3�}�C�ћ�h���z���
��5[1���g/>�7bMwT�Њ�U*\�+��&(��E[�A��K��5w�̕`47_�g�J����&��k��)48��+��K�&�����ѣΊm���(xG�}�1�I i�]��s����3z��%-�-Q��=��ۏ�rs��e�ήi�<N�����%��eB0i
��1�Y�IR������]$X+u1�'�%�i�V+E�7�E�U=���Sd���B�<4Ex�-�������i1O���_sX�~�?�Y��j����J��a�'�Ɔ�aG��K��N�j��a�yV����dU{`�Y���Q#�������������9G&$ Z�v4��	��BцL�!2��5��<�j�� �*?6��f���4v�D�n��^�]����bW���u����r�b�ɼ�n�o�
Y�Ÿ���q��c�-���J�-V�T�Sٷ5E��!
F]��P!������������E�<���YG�̪Я�9�k嫂�i9g{�J��/z��+4Q����%NvVp� >�d� P�Yw�KCj��x�X/���!g�%/� [F\Y�T��]�0�O�YŒ����k��(�WE�;�n��cK[�*��E�G!�J���̐z5�
�GҖ���4^�k�}���9/���zi�uF?���a��.�c	�����n+�}��/zC&;�b��h�5�3m��c����aQ���c{�5S�y����ܵ_��~��4����+O���W�����{��,,8���C���6a5Wbt SG_����ڑ3�+���':{���3��u헠��ܕ�;v�o�]�b������P2�#��&�F�κj�ϼZ�z�&��q�ЂK�#�F�������j�k�?�kP=�zf�͖谘UT�s�	O"���D�;�W�<��� 9�J��ݾ���3Ğ�����֥�S)8��pM��:Z&����h�����|O!�`�`T��=V��`\�P��>��JeՖ	쟴XlxV64EB    2873     8e0x���CY�9�7��6��A;���1��,(�Td��Xu�3z˲^į6���bv����Ɉ��n��T��6��������0p� ��m���s
�7 퀱D�G��>��\���y�3����%ʉ�g��(e_+��,R�<{�8�+jp"
�(�N�B`���~r"�Xc^}/G�Ln�Qc:��{�?��2�ϣ��~&-�y�d�����b4�ʩ�ߋ腦�b�!a�Vyc��O���cC+��ަA~�VE��0\�e����Ź��!����2e�Yj�� '�Mh�$���5�,w�SJQз}��5�����z?���%��D���LT��݉m�������Ј��˕V������3S,��8�-��]��m�0����0N2Y��<��$c{�;��/&ˬ�*�l�!>������;PR�_F�6�w��z|;��,/���O�d�ܧ�/x���|���J����*���v�Q-`�R�+n�B�C�����gC���- |�`V�g;�v�T���@ءx��ߵ��x��J���'n<gr�+.�)xi��!/����e}�4)�����9����P@����c�l�C~uDA]So0�蚏穨�s����.ͮxUR��0=�Bd��o�5��l����|B"���Z���[�!���l�
����6.��g9|��c���Ǘ7�$o������xp���T~�B��ӳGO-��;���i����[*�	 �u�&�>���L)�������u�A�,������bS�	����E)�eRRi�`�:��G4�N���8�ԓ��7@��	V��������l<> .W��VlC�
�v���X��3$��?�}͐���`��zm)�&<�����]�&i��t"��������2�(э�7����̳@�����k��	<�M��>!��Y%I<0�-�ȣ���H�p�23��cf���z6�JmA�(~�_����?����>�{��QN�j�W��FR-�:�<V<0ZS�)�F��m9�T����F�d��nQ��|E��Uk]GA�eu���H!�Z��hV�L�x���b�y�x�^3����Hc'n�e8�<x���!H?YO�>�*%+��q�C`��N��F��v&7>fY��|��ƽVe=*i<F�L4�TJ�.\�'�d�Y��e��U���x�k�M�j��q�2[�f��Һ8iǟ�����A
]��ZߏN��k���N4-���j�_�`d�jަ�O���.�@�m_�7�n��,�������0nP�r)�_P!*�[���ޛg���?�ˠ)�3��n����]��W��Ǭ�6����h��b3_��MoW�-�nzN��j� ������c�퐫��}���ZP�rV?��o�t	-�$���c���T��=��� n�V��ʛl����,N�i{DM�ڭ�NDB[Kڑ&=H˓&�`lPVO�j������/2�)�z;���q�o�������Adsh��>q��}ŕΊ��j�$�+�	m�+�>��_
���hȉ)�`���i�z�kz��9�ʾ��}'�X ���*��y����A����a	���}:�Ԛ���	�]�ѯ�l����	�s��shb��沮�C;P�:��B��7�d�G���.
hUr�9�._������͇dAOz�g:��SӘ>��+�4M%���N4�gZ��8w0���H��Pr9��7[���A�C>Q��|�2�p���*,ݜ!�Z�{n��+�g��sT�X~W:a�#J;����/����M@�5�VWO���舂�h7�D�	Z�h���]}C�@l�)@��0�旀�}�Z8�@U��O%�BP�����&(s�x��oA�X�ߚ8��^e��-��0�W��?R.�׭|s�9�l-�g�Qŕط��M�έ]�;/{4)�"�Rp���ۚ�F1;�=ޞ�.IL�X�8hwԱ� /o�	hAB���r����P��{�7���e��©�n���%��5��"Ej$��N�	|3OI��"�_Ag|[�	��=���3�J�-f�^��!|t�Z┆1��9V��%�("�n�^DɡԷ)�%Y�!�JA�%�q��P�y.F�_�l� y&�eG����˙�_n�-vs�B�B�qs�%���Q0�[��~���]�2�Fl%=��`@8V�ƶ�EB��&�9-~/M����u.��ٗ��sDv�?w������R�9f�G�i���g��P� �$�/7Jg�����~�/m>IԪ�