XlxV64EB    1b51     9d0����[I�Z��S�"Л��-"mnw����V�~����%��C���{���d�s8s.�-�����X/�,OyM�E���	�7�yu������QD���A`���x[���B5 Kdl�+������NT��R�] �J�KeI�_�����^�VR�&5F���/��B(�a��=P��xL����NL�
�u_�}3�V����A�=�����m�I�=R�s�K�3pyb���Ȃ0��q�u��	���%�	�AҰ�q��>j��,���b�BpD�	J�T��t��9�m�#�O%y��w��:!�m+��[E�$�QW���΀�k,J����L������Q)�s�WI�-x�k�V��,�tA��.��P�N�S����sNnxMbj�1��d+{�}���^��L!�qk���ZĴz��킶�{�ũ���z�>f��QG��S�N_�zi�G����x�A���2��6���}��"ol�δ[/G��A��P��ٓMMc�����	���e�S��X6gq��=AX�����C��'�;�i�=�ԍl�8a*�=p��~!�dk�Gx2�1�$SN��(Xk6���������׿e�Y��Ŗ�+m��㘦���\��<w��y^>Y���@W��EJh�����|"g�Hg���a���%��3�����W�tzD�4Qg�����Bd���B]u�/<�b4Hr-lzqjך���m�^�����~a���9����jy�]��6v���)��[l���w��Vr'n����{��A]��|<��|1���/�,��3u����1��^о�����P�� ��] T`g�� �3|���v� 6㠚3��P$�v��e �_NAg8���_��T��9 J�,�v%���^���~����rCf�MB�z���(�@���U�.~lm����{�Z/K
�4+�^�
�#�������70��ˎ8���h\tZZ����O1.��Yj8��(�GLܜ�>�>��I� %OҘ#F#�MgD����8hJ~���J�H	��3�� ;	�ouv�����<��|I'P!��xR��������ru[L���%�� _��g��o�-�=�j[��K�!���������=���2��)*�a�;E5�k�Gl��jñ0�)#��J4����դ�?�F��Y��r� \�%�<�u��M��Y����=���&����^ު���ؤ�-�,
�����!J�T�N&W��J/��&-����#l�.*����@��G�d���ďŝ���	�2�B[��hrW�e�P�G���k�\���ǃ�o�8�gD������0������Én�aX��2�W::�Ҹ�A�HC]��.��y���w��K u�h ����ѣQ�l}t���+Y%o2�Ad���P����n�����.����R�U���V�}�
2Q��R�1�\�%����N�`�	ƈ9G�3'�E<�P΂�ܗWd��)�a!����oF ޻�H_ۉ��7䯖IJoߠ�<z�v��;Y�T��@�t�\q��v6�o��k/b{25s��7��:{��~Q��P��1X�Ӓ\�?AshJ��푠N�>��v�����x�|	v6!��R�^t���z���ߠ�DK�KM�͘(���T���q��ii�����!����a�b�>�>��DO�����X�BHd��W�B=���jM�x���51܉!�r���*��!XQɻ
�ih�-���bzq㞀�0��@�M9{�E�.�����m���_T�l��J��Y爫U�F�v%]�4g8��ԭ%p�i0r@�_[:a�y�^���X��\�;��|��~F(���&<������0�_嫿O��b3r��~��u�`�ip�>�������چ��LX�^T{����7V2g�Gl�0\I�{����ݟjx�L@֚A%�i�.IG(0R�y��K`�`��{���fښ?�8ع���n��Gk�� ��R��H`?��F4�W]��t�>1�Ww�+��pFD�=fО|�C�5��	cƞ�K�c�A�Q3ɲ\	A�V�����;�8Y(���^�z�9(�8L�n\A6����y��W� ��'�$X���x��v
|�mH��Cn=�2:w!���M�D|H��B�f��-�n+B=G(}�!j9��P�&�O�B�B�t���鍻us�@���D:���3��*���UM��vt��i5�Z�[�J �EŞ詌{�@Q��'�s_=��ǃ6����Bs��ӵ<��`����Z�KI<^�P��ο����^�����C���O�ðZ`Z�����7��L�3POZ��]�jN��C}��k;���Pu���c��z�:���c:�M�S����S�g7������m�S���$��<%���2p����1r�	���p;��b@w�4A�7<���;�i���v��~ 