XlxV64EB    2e73     cc0��8PQ!�Ɉ�>�o*�6�1K�CL
|H�=��Ԥ��a�Ib�~d���(h}}��8���['S,��A"�ICU�s�$�dZH�3�=�n�Ų!0�_��A	��� n Eރ����N�ߔ1ȿԉ�V�j�����N�b�)��
x%��n�j�n���z=�j���0�~i\�^�1��L�.5��l5.�+� ?[B-n�B�2`+��Y�5�W]G�պ���o^�WX����rٴ��9I�wR�F"���^�h�NsԿ�J���
Dv�p�OZ^���}섄b�����j��p��[�~�E�0����}�*W��J;@���ݟ:��;w-���'��A8G��QUf�\*��`r�c�e�3��)�U�ϩȣ��S~0#�Ih����ry�UV*=��p�n ��S aSo�x����7)}���/­���@��o��HMI�P�ZC0mw4�r*���`)�BLȨ��v�ـtNG/�͙����E�O��$:�(<�z�\{5�s�zc�%d)Ų-�{�S:R��o�V���<$�k���&�P�x�Hd�PߝW�?���K�~V�Iv'F���R]:��$�� U��<7�V��Q �ki�xꊈ�X�|�|E˝�����G��-u�[�*�Y��\8��B���d铰�=��<�6 ������.1>��ȿJ/Ę�{pr�Yj�E[	��Kj�
 J�1e"�r�ڀ0pjC��fr$�p���I��s���S�^��s��w�tF��<~�DΖ�2�yy�FQwbV���T桯��F�౨$a�Ȣ�a��_ȿ��`:8�g�L��ǋ�+�X#�b$^�&�D���&1����Oc�#�m\n
���m�42)�E�wR���F�������y��4�(g	Dp�SS:��G���
V_��>�Vب�q����Xٴ�������-O�Q=ߔ�7*���X� Ġ��; �QCב��λlQ��t�x��<�O����htSq��0�e�L�7�G�+B��=g��m��O`NE���� *�=�����&t�a
��3h�� 1��:3�X63����eմ�`��C����Juu��F�kY��}���t=�R�Br��������V#��
w��K̪&���/�Ks`g]���\��O���pe�?�4�׺PX��"l���Fԍ�ͮ~ց:�lDc�5���6k���R�� �7ԩb�];<H�6� Ԗ�ULn���g�w���xd����Ԝ��
��3�eG�����Ö�#[Q)��hmd6g^��YO�[50y���ԋ������j+	��9�����u��"x���rl}G�)���ȗ�Z�+^V� f�F@W�q,���lnʂ�rI��@ߝ�z8�b����&:��%�g�-�Tl"�<�����ɝ"_vZ�*�K�4��폽�)�Va�O���t��2��h�4Vl:�A��E)Q�:����2�O!�ei�� �)���3��m��^u�����7��m @��8i������T������RwHɪ�.w�!�D[ېn�^2i��G[��FV��V��[`��*EގۈhC����MٯzS�g#�9�fB_�Uu����8;�0�\��y=�P E�I�������AZ@;���V�l2>�����(?2	6#�ޱ�j�{ 4^~Q��@��NV���)����k��� ��/���
��x���bX��aǦbY���,��ؑЗb�U��
�o�v��7�G�Y���c�iգ�*�)���Љ"u�`����Lc���g^zvl�g��Ʃ$�rC"0k&��ߜq̅2��7X�\ ��]mO��n�3�2��(��Y�Ɇ�����"w�#��� 8�K	j�Y�	}"�geU}��o@��d�.j|uq����{Vk�sO.���B:�N�þ�t�cl ���u%���r�3�ؠ�Ԧ�0޿TX`��bpG�ϒ�՘�+5��&x[�vo�4-��X+�e)~Oy�W)XH��֬� ,��q��G�d���7 )㳥��x��fv\Y_���ǲ�b'���P;��R���^�M���ٕKؗ����uN ����^�D<��F��ˎ]N>�[Ő3=��jF�|��h�t��u�T��A���Y{j;��D%$/Eid�3*x�w)9�q���0%� ��s����^�t��E$����ƍ����o�����gK�]��}hXS�`���r�i���)��t	{�y7����W�����c� �u�X͌����c����BB��&7�x@`p��vr��j��BR�h�+ O�.���R4��
�=��WbR�D��M)�AN>��5���9��5��΢�3�.�����{0v$���B��
�+u�ױz�k4������Z�G���_����ѳ�>Ŷ3�Z�����ih��QL�fF��_v��q������W�P�=�l��˪��Y(9Y��_r���Z�ߠ��JV��Z-Z�7����k�����xY^I�t=���.c�	y��/D�-�,6����<��'y�]�R���F�;B/���z`���z�ZL�O2l"=o�9?�
H���*X�.�����%v>�4�,��k2X� ��i�ұ�Xƨ��wm�����/j��09�����4B�,��	� u��C�dw^���]�ҵ���AX�gT�m,	��z�B���v��|���y�uik $S0�t/�Q9��U�n�&�TώK��pC��'P��RX��x�iT��J��ʆ������� ���$Ѐ�H�M�-�[����?�mWF��/9�Z;M��^Aa�ڡ��.��^��:z*��D�U:���9����YH3&����@�<��|g��Td!�zJ��aIk�� �4"2]XI�'#˱�l�q��k �v�e#���Ϣf���O+���?��\T৿౬�g�.5����ړ�N(Vw��j#�� h�|��%j��`��'�!���P�j��QWQ����]��S�;d��� 5&�.��ISw4WB�,
5�-��H��� N� �E�a�(w�9"�4/}�.o�1����M�eW�o�Sb��Ғׇ'<��-��	�ʃh�:��O��޾�;��P�7��pwh��3w>�F���)�Y8�/mw���{b�р|@=q,v�����ڗ �.��Q�%�u�U�[6L�oT��z��I�O�����9��·}	�4�̨�L`�Q_�����/