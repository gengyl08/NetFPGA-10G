XlxV64EB    a70d    1bd0�NzQ�U-���`ϛK՜u����?���N��.�F���Z��C[x��~�/[��U~��xm������F-�T�S�@'��x��Tzb_˖g݂C��+�{�,&Cf��!sOщ� �6w���3<#5p2*��p�-J aD�t��37�`�K�"�-�Fl�ܠ����8㲬+�U"_I��u� _���,HΓ�}i��X���n^�a�7Z�r��K�S��1�O���d�e�W�V��d\�M/3A�Í�j?���S�1.���͍x�q��lÛկ�S��a��WBގ8r�օO(N ً�YpHJ��Sm�|���+q�]���7I{$@��e�x�B��=�`E>�601�����C��ΊI�4<�~W<
�Ϸ�~��8��W���=tU�c�mvwI6@ײ/������,��xg8����I�A��`�9��deǏ���w��F�V�h�2!P7-פ�
(G7�#u���~��5$�~�{�8���^�����y����B�X�i�HP��+q��Ç�����^��\�b�*����4b�nX �]��������<LT�T�����EX��Z���s�&x}��dA�_��9�Y�a%jpI4���U��ô�/��|��d/_�L�ۺW�����i d�t2�	8�2�̳��$^"�D�p�bE��L���8�1���l	k�Υz@������v;���B�&�9PD�>���Ee6�H�h��A��X��E.���U)>�jd�6@qz(�Hx� 
���xc��$�9T�g,�Ie.���t����@�0_ѝ4u��I��K����Tv-x�j�$^�G۽�W�`���칼��c�$���7��k
�\e����פ� �5tB���FR�(�L�S�$>��kI^��n�11�����xG���i�D���4*����S����YH^,�rV�E�Q-�h�>������?R ����i�y֖������]#��12	�f��/s�˰a|��S6E��!�4$b3we`Hz��5�J���L��:D��na�g˩kw����ԸhV��8+Z���"�~@i�X�4�(Q�.^;v��q�>��7�-�h�s�0��0���),p9�8�T3>��a�A�f��N�,�"�����h���t :c|.��Q�� �v�!�q|"���?a�Gv�0wh�|Tt �^���B��PBp���J{��B�U�\�3��9�tw��0L�� � <���>�]�+�,�L>&z��t��g�"���dt6Ϗ���F��N{sy3� ���/+�$y}���Vz���!�e,u�n���c֙)�k.d�Y�қ�L��oU��	�S����K�#��"��bQk�o�	+k����7�d���.
_T}.I��_fJ�$�lB�n��K����v-"��������RO�r}"�ϳ�a�X��HDn�	��%5��Ot�9�*i��▤7jL'���,S8��y'�p\���i��K���`��e��^:0ٱ�HZ��,	*T���y�k��Ӗ��:�F�� �d�^��2ųNm�X��s���m��bmi�7�R�G�L��V���9R�B�Y��gA٘:�A�:ut�u,F��N��Q�.H�1VC�$��F���jj��b����g���).k��4��.���([!��_��#��uGy�!7�t�;��u��#d�o%_]=��A��K/�5����x������h��v���}�B�)�x1fJ'-qGmQ��3��󽛠#���UsGI�N�#����z�H��ӑ:�>�'+�]&�ԨX#I�؈���%�3��n��V=���B��w*A�6���w���5ȗ�˳�gC���V�5<S�H�����0�PX�01�f�����g������=���t����
��h�%���yQK����@��Bi��XSZ��~�6���ˀ0bpw�<1i��k�_hq~Y�'�?
�s�iK5�ŞF�,$^4Zk�Ai�{	�\"/���]����ʳ_�&���)��|�خUZ���CP���.��o��Z���>kY�
MH��4�"��J�6�[����&�o�{;��<$<�bHWm��Y@GP}�Z��,�4�Q�#z!!	v�����S��;-
���EW�(�g7C-��
 $�js1y��� ��*�Qz���J���V)��:�@@#Qy�2��,]��ҿ��^QF�"��bD��:ƿ���K$��X��aU�"��r���=�?c�ޘ�Cy��=vs�K��K�(���\����e�OB�����]�)����m�&?=(��Rf$��Zf��4��ձ��9#m"��ߟ�
A�n,~1U�|�7k�A�&)n@u��}"Gy���2{�QwTuY?�!D��)�������܋��1�:4|9
�̿y��h���?xʹ����7Nx�\��Q>6~s�#���34缢
���I~����9��I�JP�� �QfC��d\�[�H�)~�[5/����n7u�u���F/t�7��K>�힎���`�<߭����^!3�@u�뻀z����˭��z���\U��eq�\�-����;"$H�̿ȡ �E��$�גU��y��))��L�{]3+l�XЇ�m�Ư���>�̓V4���:���2b�p���@�����RG�H�ŋC�\;���I1�:L�v�i��
b�[ '��1��̧(�j�����6�� o�X8�{eP�Y<�U��+���HԢX~ܐ�1{�9���u��"VӔ���T�ܔWa��:��3��g2�!e�j����PB%�������!��+��v�ۍ�٘����f0Ú�+ɦ��}�/
��("��R�'t��AA�Jٵ��M`)�u����_�Av0[0j���Xm�w�./L��m�j��.ris����+u���b%^14+�h��l�����E��T�?:ǺX�(_�I���o�+�q�w��J��~�Y�7���<3E<�VؗEFP�e&sJ��L8��șډ�:U���/��>`v���4�DO�S�A�S`�_�d�\�vs�����#bN��#CH��U+%[3��	��c�*3N�va�O���6z�,\i�}$�-�JI�s~ѽ�L<?��V@&-3�ӉE�AzӧB�t�a���+�=�]���0��A]��Q<�`��^C} ,ѭ�(�6����<^�ܩ���2rWip_o�։|t}�3�̙�_��{�J���5J2���zw}�A�,t�N�z)�� y��j��qr������_R���`���闰��y���(IwY��Nv�Ix ��n&Q�V���Ǚ��O��-��BGT����v��,ȇ�fX��ę
z����H@����ȿl+0L�I����ӳ�<R��n3�z���&s�Xs���;��L	j����g��0���s�,�cK&q�ny��AW�d��K����I�ٛزg
$�i�|aD�
�0z���yK�#My�:��O"`����3�}�bezD�bw Eի��s�d#�%��8��J{轂R�0˪��D
y|�4^}o��)�2R}֦9�\֦ޑg�	7y&CG6�1�!�ZS⬅�у0�7l`�i�8_$dX�:��U,-�E�-,>�f���#*@�#���O���ŭaS�1�������D����b��߫CG�����=Ĉs-�y��*�,3��r������a�2VP[[hH	��m7^U�X�}	!�ogW��\w{ `�&�_R��Er&�+Dr�p�ڥ�s�@D�k�4���B���t��mj�t�=Bt^H������=�h^��!]<g���bԎ��St�x#[T�icG�a�K��q��|{HbMq�b);p�']玭5be����!jૡ��B�#�G���$���{b9�:�Vr��X��|���B���Ȏ:�J�-V�`Jy����\�A;�`nw���J�Eⵒ��:G�(�7���
N5H�fA����� �@qؿ�M�	9m/ۀ-��G���!?(���a�<>.����>]l�t�֧�]��Nӯ��T)�Ǌ���˶�bDZ
�j/0�e��+~-�{XD�8��h5W����C��Z�d�8���6X/n�H�z9*A���`d��^ZR���Vw���$�->�gu6�F��n�`�ى*Cs��5lL�0�CB~E�tV��%f%��T�i�
�{�$���eX7��d��M���^;�8n�#�����&g�eWɇ�W�Z	����A�R��ʇ\j�$�����$Mv�h {����zw��I������p��`���f��;�vZ� �0�X%U ��Y�L͐FOҞR�!N�uF�[���j1�h���
p��
9�'����#\G�fkt�g\Fߟ�>(-w���S�j�I_m����(�g����Ƚ>������}ȌYIв��!C{�UY�;��s��\!(��o�~��1��7�����؟O�䢡/DL?	 �\���T�I�v��O���{k��������R����!!��`�α�G�\�{�59B�����0G"�9��KI�"�a�[�.�@c"H�r����d{l� �ɥ�hC��.�h�?����r�yb]�^nRR�b�j�|��6��_(ր��&� ��C(�ck@@|a<^��ܹ�e�D#�]!���)4�O)�f`µ����=����+��"�[�:�%W��p��)�e�W��w��o�x�`�� FV.�0���>���e�#c����hY�!w+���/���uq?̘17A��H?�>����&Fv��9���S0V!^�;Q���c�>�};lX�U83(�n�[ٽbaԄ<d���b����sZ7�up��V�~�R���joy���gFK���R��{e�=J����׽�h?ψ^������Lo(����-c����E�(��8δi <�L��3E�eB�I��jZ�¤���ˍ�3USg �G�1�2*��Qۑڷ� �Z��u�Z%'z��E 8^�FZ�sgŎ_"�B�u��\��T+g��D�U��r��π+�6�ދ������^��. ��'Vh����}�&�c�R�z.4�۔8�`4�̊``��	�'׮f`,�'1@�7���@����� W�;P9���+�(ڬK��'@} ,�l$�3���0I^�����=�b�ȥ��ދ?d�]����iP�[^�E� ��3�5��e܊�c���X}=�Ld$�|�o����vO��uĦ��ù
2�<D/u_
w��㲭R���ü|;����+]��o�:�	a?���T�vp����B�i�����;o�<� �s�$������|=��p9s��Z�{�I7��I��O�8	��,���z%�ԙ��I#��W������Є�X��qH��r$7���J�F�m���×L2U,�W~^���9w=W�]����2&���ZY}R6�ю�� �ĸDZJFqf�����Kh0�?�w�c�1ѧtr�
e���4`:�z� T��(�)�(n�#3�K�Uӄ�DGE�hj4)�[n�� ��l]��ܕsU�[��⏚��?�#�-5>Ш��a������ZÁ`;��I���q�������R�n'vzt`AvW��z�F�+�-���Z��9�OQ���=A�z$�a����;�Ɂpb併?���������&\�TRP����\]u>�n����\�t�<���ݗc�_+�j��u:9F�3:}A�6�6��]�Jp��Ifеm�jh�/�����_��53`�9ꗮ�B���mpf߾u����B�1��=WR�\�!e��Y��'��҈lȞ1��&��7r'��&��{���}�����-����JW�t�妍�Jͮ��+!t$�Eݹ�Ds��鲐9V��Ӊ��lh�>�sf*��x�G�E�)�˓�V�����G�l�w�/%P]��c�W�%ଐ�q}R$�k�r��W�]�c�?��^2�4��v	�'���.+��
�X% bI�&lP��.���n_od5o�D���{��!AC�Z��HL���&PŪ'��OJ��\۔��,\,Nq{�NȪ��5
2� �`W���p���x��,�^�m��ktz�{U���*$�����9��|�EZ~oD��A�>�j�����[�� K�i�������h��r�N���2zf��Z�Oq��@�eo%3��p��\�}}?����Җ��R���G��������K0��]"�0ܽ���(���3�|���$/���^��y3��$z�}��m��E|�f�\���,���/A*�3C��9�ݻ�S�j� �N��um����.�%��fܿzE ���]U~��aWn[��7Ǵ�}X0WAd�:�y�ס[fT]���{h�~�+�Wđ����%�b%T�(�]M ���\��K����O��X<]�ğ�EFq��J�R�	�t0"q9�B��g�Y��!��8p^���\5�����%ih�̸��Q<��ђ0D2�/��4�zp>դ��]��^�l���^�TӀ��K86������hTze�o��)鞌G�P����
�M�&�I�!��X�1䖑�����ʹSUu�!5Y��A��v]fSSE�= |<��Eޓ���S�(�����?��%gy�hO����D�E����9�{�M�&��Ӂqĕ
#ʭ�@�DU�y��CƵ��>,�'4��J�u�'JLf���/A�v�"�R��ҩUk%�C��E<� ''i�P�L�����Z�N]{NZ~����si��kle	b���E2�����?2o�+.�����Ŋ�5�)�.0͵$��@� �'�&�:읤Ќ�nѻ�&�H�a����\�	�,P�1�JG��k��ݑ8��#Mc�6�K�*��;�*�ܤcG�p�t�V������*&J��+��
+��Ko�"��,w��r[3n��n#��Ǝ)�h�cG��
y���5�3��h��0u��;����g�cA�x�W����u�w��(����v��煓τw�K