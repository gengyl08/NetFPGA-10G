XlxV64EB    fa00    2ec0����XqI�.�9���j�ʃ����̻���L~�_8�����h�)�>��yg\����}�M�Pq�X��,'�#4���W��|��3O@2��2)^m�@�[�m7����0�KO��7F�M1;y�`I�,Q�
��WL3;�0�ro4O��� �*��}z�e�I�u�F���'���K²�hH��]��0ޫ�t��'�N^��4apެ	�+h9.�D"�������pI�ϡ1����8[U��ה�*Ձ�[�6/��e�Lu� ��X�g�E�+�8Y���n��i�%-�[zL��_�bmH�8	�I��U��iw�������h�WN7�~��(��١�]�	�KW�,����?M��	{��PHY�荹F���7�Il{�CQ�Z6�����|�6%X�;e2Le�)��'1n����kS`�f)^��Oɀ/��S:��J���.�l�/*�)���G���`;u�^�QY�>B��Y)�X�[�Q"���X8��V:7�`����Iqx	9�tM+ȋ3��^���a��x#_Xt����j�-�RO���v(˫G�}8����&�4��@Utг��{kC�1��gґ�5�V7.>S�T^5r	u>�kuY�s�th��-�'s&F�在1���^_/��EK���Sj��O�,"!�+��b^���9�T�� �p���y<r<jnG�<=�~����au���2��9��@2o�����gs^Qx]�Ă�G��<.���Pw�Y�|�a�t!EGb,����V��D�WL����$���z!��P�UW�f���!,�tûeM�Brr�����_��J���/v?4�W+h	򢠩���t܅QM�\uƌ�t�?��������a"�I����K�	/V�*L:��.��q�x>[A����B��4�z������`�ڶ�|dhmW�w�����c/�M����8�&�f�Y�`�X,���*�2p�Bz���ԋs´٭��X_������U�5%;��_�8�eG�ʺ%Й��+�[��:����r�(�s���vyKJʛ�-l��C�:Pp:�9�/��3<�B��ϴ�x8n���3|�����j|�d��a�or��!�ݝ�aV�� �Pm/!�ٝU~!�p�Y��Jqu��@�i�׉�^$j	�l�(v��в��/�@��� ��-�����.��O۪�(� �y�<�q��i����4"Z����D?!L�%:<"�7[��]����|唼k+���T��g�s��J8���3Ҷ��w̰ڀJS����i�s�m���7�w�N]k�y���+��R5څ_$��-�!�V��*'C��������ssu���:;[m�(����8����#��sМGǌѬ�����.s<�?�ȏ5y�n�aA5Z�R�Z[Z˚WԨ���k%�Zt��^'rO���S�.d���²d��4�~+��?v?,��9E��E!�Ӹ��N{h�݅b�c�+4�G�q��I<�m���v�x|�����"�y++�4�L��>�`��c��s�����/��6�8�V;u��s�������f���m���F�^���A�r����s;7�0֤
݋D�9,/9F��TB|Y�#4G�h�o�����q�g�'�`9C��o�gm�0�L�g��Wvݲ?&��i֍��v^7ŠmiPQ�rMJ�[Gg��G�Gs���-������G.�������!o~[/��4��4�z�VB���>*
%�a_��qb;�K��;����JvMl��<9��8 �}X���?k�Nl�/�G^�/��0&��N_�$�X3�����N�G\��<]�8��a+����v�s�oo��O�p3 )��i/��_���ș��=�4_l�[�'��U.��Ǐ|{��"\������)�&0zL�a4���a�6\�������1.��IZ���^h��5��T��*��������XLC�U�jƌw7܀�Q�h�4��0r+j���0�v�QxC�<�PR,��V6e)�H��^	bw�d�0�h��^^���>����UC��a�/��V�mЄ������WqP�DCĜ	R��1|�aA�1�e�=��X~1K���#UM�>�8p�}ް��>�霈t#G��k������k3�W;���	���6 V|6��6VO��LK� ���*$��D��e�2�*C"�����q
_,�-%���xQA=�s����&�<��k=�@��eE����NE��b�}�y�{'�-_&:�9��Qhdg�����;&=L.˄�z�=�)���K_}'#ޯ���tMo�"�����|��I'*�"��/V��k���T�4���2����ɭ;�})���=ζ@y�Ũ�^��D�+.bD�%�h�幛U �|g���X}m�ͳ�ߙ����VZ�VS;����;�{�9bz8k�U��}�Ga�%+zw�v��}���7��n���w<,����f*�Z�bO�դ��.�����q�m�<�6U�X&YL3��</"@3� �B���yr��[������4;���U���G���.�'R�kE)���g�rX
� %�Z�*]��UK�S<����.�!fl�:Z�Z�e���l�"b�KnXQ��]��s�fM��}Q���Uv�6<���a��{7�V�	��:U�����Օ��-� n�->| "gҍ�)0
�N���U����=A�M��a�Y��i�vK1��$��-o���[� m(r�H�Ҟ���(��b��;3[��#\��(���Y����'�x���͜;"�Ƅ7m�z�Յ���Q��pcZӃ�ض:�'������B~�&E��ڥW�-�&Z,�5�K��<`���&b�ly�����6g��B+�6-��p;n�:|���$�У��~�$<�ti
#����-�2"eE��`�v��r��V�U���i�b��e�Ѡ���MO���{�Q(�5�����M��Gv�{/�;7��ٚXl�T�~<@R�Y}�Aom��ӝt�>����ʕL�cY�`]����,:aUN������ru�������{&���8^�G�:��� [Q՜rpaj���X��o���2p�x�=k�G�OEZ�,��Q��83�nI[d������r�;� ��[ |�3֍�d;a�8�KL��Uc�Ib�Nq�"���w��`�lQs�;Z�I����qbpA=5oVg���$e���s;�+)[��R���rp�Uf�\п"�^bV�p���!�C���R\ف#��4v�:��"����U�����&{.����U5��p�� �#�o4d@�a��=컊M�ѭd-1�����w^p�-JGEV�������*:�6m)k[�s9Ps[�tS>����#�JD��B�c�J]�Q�����C�y �$���<sަҜ�
+[>E�1s2&
O%�G1?��'��s�ޜN*]]ZN�Fe�f�w"h��~�}�3]hh�{/�	k�ޓ�8>/�m
���8�7rG����LIԍ�11V·����`�Әʔ�ZD��ߺ6����jDɁ}&\[��=���W�,�o|@�Q��T) r ���-�0L���'�]�x]N�Gz�4X{��$����$ ��>Z���u�H�|�������j��F�f�W/�-7�&8��g5x.�Z��$u���Y<r��DUv��U��:�JHp���`(��������k+�l���7���;ؗ����<�V����M)����wn��J% eS�{8��o�>�;��)�T"�t��(H���OW�k����"(G�p?�E7H8�:�3��i�%�S#3"�_��E�Ī4:�'&�_��&w��E+�U��B�5L��+f��$�� ��ڳVp�9��\�@#�_��7�
�X=�,��g�+��4�V�������GcgJ�L@�QA���		�R���R�� �e���j�B�����;��H�:�5�u���8�^�[��=�MO��N�Z��gn\פJ��^�ܣ5�����Ņ G�o�q?^��y^X��&�/��̈��<��stZUn�p4;����}�*ن��z��̗���ǢYK�38��rU����IK~�Հ?F%�V��ֳ<7A�`l�Q:k��OA����ce(��H��S�����/��#��8$�r���3q 	zٛ�=r^��n�� ��p��΋�����U+���:|���7����i�������"� �c�����h��4�r �OCMZ���Ն�G�`���Ǻe���B��Tz�MZ�A|с���~7�>6&��+M���b�Q�'�6���=�s��c���0k����M�����!�x:ZA�M�4���"��h�j�ӊ�`A�"e<����-�ƈPTY�d�q��=�q�H^�����΀�.C(���b��S��NObJ������'���}G�t����Q���q���ȼ�0� 7���7�(\��h�d��=z�Gxc�~)e��#ɻqd��;�h$��ݔE-�� s���{��_�Ϗ6�t6�ȧ�X�^� Q�͍�����Al��Ԝ�A��^����{Ӛ�^�uV���.�$bJ�PJJL��~�kK�d�bФnb��D�I��2�h�QTH��ci������l��b�i�)1�^5�j���Kt4�]�0��w�-'.������X���:�p���8&i5��u�������^3f�n��^f�$�o�&�u�!�þ̗ �=�.�N�ߋ������q�K=3���j�PX8+V��[�5z�ɱ^ۮ0��C=X
�� B���&�^t�K���w��)yQ^ZLب��F���P��6��q�Il{N���k��\O����W���G�ؘO��S-.^"g*���v�2uqQ�z���)@Q���qo4+x��s���<i�P�+E(}T��|����{B~�N�!�ʤ�k�90">��f�Y
\�]��+���0�<8�l�]&t4�@)��~k-��׏�&��>Y�r)֑��1����s�
uŊDjmX}��g84EQJ�2}���Z���Zd��p�hF������B]�̓��|���M�e���Hg)
�ڄ�m�Y�
4W<.��\�6�7<^�/��v�E��I}D�i\Z>ѯ�����mL!��fo�G�}|��`[����.Y���K�2yB��x�\���:dЖ�v]i���FN�$Vm���?kܒ�sf�S9�˼�G��+���#�ͷ�`�,?�K+�����c����)�4i��n�V���q���+<���_��]�nCg�f��:G,���/D
_X��9����1Ԥ�qEOiƵy��g9�I�mV���uAL�(F����)uSo��llG�z�=�0�ݓJ���Δ<��,se2�T��b����C��a��#��,STl�WvK��	)~E��i|^T�A��J
�]ᝧP*�;!����;D��9��2㟶Q�dU��A^�H�f�<���E`�������9g�(�";�|��j���F����ͮB��,�r��;�)�kC#q���8(���::��V1� ��O�{�$�V�N:R������Lv�{� !�{�$I��r:�ϟ0$��6���`ѧ��s��������r�d�)���Y.�g_�F^f�c���X��Q�$Ua#_��L�e�-���E�SP�l�My�B��4���*�֐�J��ϋ��o���s�eֈ،��FY�d;;
ϡ�/[@���/��]-W%�a������bT� �*�*�� ��5�{�Fc���aj=��F��`�d-ϽS��⽺4ɷs�*O��R��	����?5�0�dc�O����6 Y�ٗ�{C����>����L����?;T����I}=Ce��TQ���aC�{f�ʣ�9+�B���y��kL��&�%�v�������Z�y����ٻ��S�9#z�+��_���:}Nk�e�.:��7�
�J"Մ8evEaVhu�jG>���y��p��$��`*zg�%[���#�4S�A쾖n�_#+ڗ���h�﵈n���zF3tm�#U�~!h�����m[7�����t�݃�_���R0l�����?�&/4�m��y�
�a�WU���X����QʥOw:u-�R�T}�X�O���+�����f�r�6E�>��O#�(`)�9in��l��P�C�Z����r��p�j�z�w>���`W�J��k��r���nq�`��
��&'�RĜPvCc���(Yhv\�vk�N�"<r��`�E�@an�Jx+i&=%;�Ba�"�3XiI�U��BnbD��Ge��c\!�6���|z2>I�_c,����sr�.�����U�y�?�*c��P�Njf9:p�Z�����BՄU�S	ăb��N��Z'菗vЋ�
�z�1�+���
A�xˤ�M�p�S�`%v6-�x5�Q�\ox`�-�P��I��YXu�W�]��8׆�!uT�7��o��:f�[$E�e� ��S��o�[���!����MRt$g�i��5�T�?bԀ�k����Ym!\n�T��)-�8�ĳ*��V㙶���,���ߑf�/�o�L!7#7h%CƆ��2C?���*����0���<P����������>�Hz��*�����`�;�~y��w`4�cs�����nZ�c��o�Ǭ�)��M?@g��]@	Mj�*r���)��wF�em�@�;"viƴ�ps��I��$�5����������]u]/F���G����E��I
�%T8���8��D bKa�-4G���y���hMƍR��>:HQ��?�0���O!Гr+�>��9�6��R��M�]��oއζiu/�یڱG��ZĢ&���a+�P1;�j�+Q>����(f���{�"�l/�{%o|(ʹ�+/�qم�xY>IVqy�vuK����u���4ʅ�0N#�E$����-��/�1�d���}�����&�u�>����ۙ�>zC#��ql\���I�"�[�і/���k'���>w�nk%�\�9y�e��O-�H��W�a��j������r�����ze)�qE��ⵠ��hG��X�l�X�8
�'g�z]=�θ-�ŗ����'b��̽D@F.�v�f<e,��+*�?_Ja[�$�p�K2b�+L�ח��mW�0���Ye�Q��.����
A�ٳ@gk�cu���	W�K.�����k��;��[����u�P��`S���fM���I��C&���[��rT���2������p�No{5������V	�xT� %.���*r��󵝌E��)�c"P�N���)t�_��ۈ�p������g��˺����2.�@��������%S��fv��~���&Wh��8���h�U��em�d�8R؏I;���L2����ڄ���\��|�!�
�|/��zw�Aj����4$�k���߈g�H9>���e�M`(�KnL K���$$��������� Zvŏ(����G��5��)����{j
H�1�z>�ʥ}��U�,&ASa��wbk�\Ptu�]���4�z�<���%��@�wg�0g�HX�1�Q>�+u���α�S9�i�j��v���� O-�"��;�Cy����t
 R9�kB�Zכ�cz�1�O�~�y�z�l��m*���rZ�0����:g�s�9_��ׇg���������QO�&����ǹ�{��,x�z?�K�����狂�U�6?_��e��31䓍�`ӧ�1zas��7O����g�'�{w\��Q�+�z��Rx�.����Wt������s�w3[���� a�|"d���g7
�%�DP~��L���8Ti|����W�(�u��Ļ��X[0Q<���6�x�@z��j)��#�K{�羏��M����gF�"���˷��Y�ޣ�j��/X)uh�yl`�D�͒.�Q��sԃ�m�1)���~q�2���2����Q����H\G����N��<+M7,�W3���_ҼcdtD1�%��s��h�I���]��a2�?�rfo
~�]Q^R��|�{�W#���9�>�-^񇴽������<Zxm��P��>ȑe�=a%���4*��������F>,�K����	~�|�b[s>���Z*v�h�š��6]|��h6�$: t�[³����9Y�h���")b&���[�ͳנ�����j��#������Im��gi�)���j=����^M��eaX�����_�h���܁��/[~~���v?���d�q�X�Lſ]����3?���MY7�z���E���rTE�q�2��B�`�>2ɐ���_�:8��l&���5��k�xW�/C���+' AA��s�*�.aB��Cl�`�����5��o��ek�h�vx�aD�>���0ΠF���Xس-�d���F�uZ����8�e�Y`�����W7k����r[��/��5Q5�BÒ�sdh�U���lG;}.m��gj���9�*|߅AU��k�r��I\��U�Y��ߥ�Ө~���7����0��bנ�&���[ECOdW�X; �%���測�;T@n>��j��8��A�� �B�����%����vj��"&Vkc��f򄆑!�*Yxkp}�]�K�gk�S|�҈�?x$Y�ǅy��9��y���D��WQ��۾�2o=��o��+[dV���J_�Av��~��d�X�4ʷ��uh-�9�y/7�� ��;]����2�����G�X�B���_����w�㱔 �����a]��j���uiY��tO��7C�$��?`l��P��`O�f�����(5������S��@=�����q�uf��΁HM�_�t>� ���:�T$�t9
��G�yr刮��D�FP]�!�x�Gä|i�S��$�;0.��N�V�wi�� ���[
8 pKvu��X%Ø>�n19�˺�����}n�������&�ܐm0�Z�F6n��?�c<nUe���pa�=f�辖�^?(�:o��.B�(�ij����~���5��E:mn7��ؗ�m��v��@'=��I���Ĕ8"w���44�s�9el�p*�/j!�##��x=�S��Ia��Ќ-@���ln��d���w��3@JbqY4Ǆݹ濿����\s�"�����@�]��+�L�䭷j8����608���I�f9uc����඙E�+��O��\s���a��}^-!Ⱥ��Br�E�5��!����=���uӏ��{�4��e,���1�~VE.�� ����عi��I�"��M�/&����c��շT<6��_%涛��}`,��G�F����n���V�r*`M/���p�м������B�K�v��WA��C5��M�sb�<�G���?�@e�y�{�\ v�n`�|�]]����KO� !��Zf����"�{�W�c��ty+X�(ɼ�R-{x������ê�ե!�������m��/�58kb��m��1���ʕ	���O� �@q�?9�r�v nP݈*��V�!�	�����p����x`
u��zn;}��Z��Ȉ��OGc�cc�If��,�dW|Kx������:�3QN��_@��`�jӾ������ۣ��ar�}��
{ea�p��?�+z$���{S�ܻ��>��p)���	�)E�f\���#����5�Nv���;��`x��`Lh:,=�ܹ��p(���>����##����$�ԏ�{W�G�?��	�l:Ø�\�� �,�g1�~���Ö��g��5��|±��H6;s�ϲ}�9��.�v �g߱9���QQ>Gٹ�?s��;��8˵f�"����_��1W�zQ��g p�����;{�M�1Zp�'�=)I�BrB�����!]���������;?[�WdRy�U2��K��$T�E%Qɚ��H� � ��uU*��G�}�]<w�Q�����30�(#����FG^�vd����������7�*|�`�P]@���q�N�~J�Hl�[��s���z�n��l�����
�%8ю�P^3��[h�<�>����X���;ޜ�kNF�Dt�is��Y���6�cu��ߓr��Fn�����B�1���hv>�ս�ȌvS.��[S��	{��A�����Z���]�,F�,�D�g��|
��yd�C�ĵI�bQ�4�ZŤ�Ym(�^z�
k�Ӵ�}��]	��������3� ��]a氵��OO��$�s?n�8��+��c���� ���n�=H�o��Z];0_��q�#�O%wEBP?���d�����jB�,�I�^e�ߨ�I�G����%��)��;����p��7R_~t|B��ʅL�e�w�����hԂ2#�tG"A����
;�J�d>pD�l\�9-a�
��\��
�����S�pK�|:G
� x&�mNa�������2�>eH>�����9̖25Ɲ5��U�J�4�T��Ao��������DM��j�ɣ����nR�ghQ��6{��G��Z��]��Y��Gd"��Gn��w�g��pY�[��Z��:�Ͻ�;��M���v��drozH>3�3i��>[�N��j(d]\����i�=���m��&���m���Mu	w4E�},���A���e��e����o�C	���
�(�A?(�*����~ �N�Â[Y�
rε/H8��5]�	}�X���M��N9����KSp,���BK�LE2��V˪�C�0��
���}8��xb�2aK���n��Սm�6\#S0��%#pR��쳓$�-�fK$\�քԷ����r��S���2��r��҉w`������vvkf@�g����T�1�C����c �C��,�HE��p��;�ra��N�Y�~9�����V��X�7�E�"��´����)�q,�3��s����Y�HycR���:�Sk�O�$b/��Y����A� ���p�6A�ޝ-�_�����
h�� �0��1:��ϙ�݀��L�qo��6|h��Er�{"�7L3Z{��>{���P����q)Y��q�����/l*U�٭r�m(j �i�$ÌV��m�Nh���1��>kn�����
�+�'��^a�JΎ&�B�-�K(� �*q�?]��;c��y�[�%r�����͖��h�����kH�NI�Å�(s�\�Ia2h#(�{�on/AD'M&������������^7�]���/<��V~_P��e��r�Ȕ"�s�P��v��������A҅�j���aµn�}��;^���q��7�8<C��p�1�5kBw�e�ș��'����g���{����<:Z��8��$�Ѿ��|_t(l��i"�Ϊ&�:���@n��m���4��#'{mp��w�Zcx�-+SQ��Q�O���b�����Bp���`.�Ro�7'�bJV�mq��cU'�7�D�wN�-@O�)���]�I.)�������rU[ps�_O1�ӠS�L��e� ��
U+�?��q(d��&K�ay�]_U<�����OC�|�Ӯ	>4��Yg�JK+�#W� �=�zOvR�:���ܳ��7Ѽ��)�4�pAue�����$_՝|�\��6�w�aI�;`"%g]�hvM��	��NK~��Ph-�Ck�JѸ���S��>p�r� D�p�v����~�����eK:Dx�ݝ�f���v<,[�B |�� k����y�@O<l���Ss�Av�8�*�(��^���F{v��P&�9:�0~�6�d3Y궇u�����d���x�h���O��{�N���T��XlxV64EB    63aa    1070�U��	]	<�\h�:�$�%P|�5\G'�l0��û��)g( %fi�`�ەj1q�J�ʅ��\����W�ƾ{�#�9xg;��)5N)�E���9'�eӞ"3�������WV��i�0^A�����<u�R��K��c
(���GҶz�Qb�y����d��a��9{+j�� j_p��{e��1_�}�=�*!�X���?;�
��W���*6d���u���^:�b�ò$�/�N������z����;e $�t�E�7;^:�(��S���L��K�� _
͖��7�}��66��a����f+=��(�8ᆑ��]Gt-��o{El�t{�����E�<Ѹl�sU����e%����:�!ϣ�U������j" J`��4��4�6���,'	U�H�W�"���$&���	���%���^6D,� ������fV�]�M�3�qd5�d��+�<><d���%б"��s{�o���Қ��H��R!Z �ZV�>?�x-XB�V������i��w���C���c���^���B��W8.�Jta�`ڇ�Yl�߽#�I��/�L��\D�H8��K��R_��C��Y$�8J�q�<���WL�P�V �p��}q
��Y��T��V}&� �1�F�|��"6ʷ)�B�;:��r�ھ>�	y��a��D}�\����=֘֘9�q�\��v.�	]��-�C��R�B���|�&-k�j�>�Y��.�1Ϫ����H�;��a$3�H��_z��E��H�S�%@DEX~soeO.��j��C��B'�M��: C�Q��81v�Ϛ��ފج�8]P�£Zm��Vp��O[�h�X�L�8Q��+k:��u�,��� ���k5������͋t��q���e)�7=$�LU=q3�4�s��(��c��; �x����sRWf� =sp�Z`;"2� �Ѧ��c�>w�t�6:�lg�i3zzj�zZ���9� a"I��D��+��=�Qg$�(rvq��:a:�������!r�2�[bo;�������O��czk'	[��#;�r������_G5C8���
�f��JR�?[9�Hv⷟���0���qa)H�+r�<uA���L��Y������!���e�)��WL	�ZB�
\�k(E�	� ~a6u���T!K-��/&��=7M�.��j;�NZ�	��h9�T���'������)Ѫh���PV�@`ٝ�kuǑ���)'�-ڳ���Y˲ Zr>�è��[c�v�W�(�6��%�;��]?��X-9M�6���~u`��jg3x%=�V>�Ҕ���?�v|N]����{�����mH*��gqbGChM�}��yŞ�H������924�G�"(�;�~�y��u��Og�d�	B���Oi��+�����&�����Eۀ����YKT���-g0�KՖ0-�~�dI�ma�t�2An�!H�`~����^mv�ܽ��s�eB���r��H[N\��b|8�S��ڲ�(`o35	j���l<m��4��ψ�h�����)jA@%�O�խ]/*���KD!� �����:������ý��PH[���5�_'� �+�-�!�<�ֈ��4��z�R
M&���x7�����i`���]����Φ�[�A�Ko���Ld�:vb[�}��kðh�BΣ�u���@��;���ɍ��� ��+�O�g�����	bo�Z��b��Vy�8�������ac�����G���o�V6�.��9�f����"� ڴ�	���F亱�6����-�Ǚ�M�Uջ���>2�3#nB�7Pd��қ�������Wc���|z�^�K�
�܂��Պ��v\�SJ;<0P��FTH4s��Z��,r��l�Lv�YbG��W;��
�NFG��r��X�4�i��T�&��
��fI��~���Aj���]G�2��A&��p�9��9 Z9�¬�1���iL��e�n�Z��HV�Z��7;��R#�zH_[�z@gX�1���@p5�q������!�^SK0���k�;��T3t����z���	�-����K�Nt���7�� 7e�
y���?��P`���t�'�f��y��믌�}�x�)*/�[i#�t�����p��.҇z%�GAqIp�}#eo��x.a�p��`�`�`��i���-�}��[-,��{"u���p���q������]��q���,'Y��n��1X��YD
���z���WהGo���M(A��X�$�.�v�s���n��
V.^�م=��2+��SқU��4 ]b�>o�G�������L:MՁ
mk���u�l�����q��_/.~�`�ɂ>c��h��?ܴ���Pvr�YT�,�W-��`0�v���bK���1cNV���=�D_�&���WWU>8����D�C,Z=1��6:�v'��� ��a��y�=�:a�h�D%'�9| eI�sF�c��aڭ:�x��5���p�UoAj9�H��z;�K�<M�}������������ۯy ڥ����tQ���Sm�F�����)"�w���m�j�Z��`V�U�H�
:<�Ԫ���X*��z.(Śc��Fv���y��*�y��|/?��/�6��������R�-o p�x��J�L�lX����`ݤ�x��L�;޲b���P֢��X@Zk���p���=t-�hr�:ŷ�-���s,�O��3�ǫ�Y沯"��ya�럋�3J�198`�r'<��ͥA�K��C�@��mz��e�i��4��CI�9��Jqz/��8���fƼy*�M\��%���:�ă� ���Ep�S�V�h@5d�SukY��E`}(��>��)��7,�8��b:����I���ѹ�f�Or� n�C��n1����m�$�)27��CF[,����=҂ʁ��brǔMFU�@�yY��Yn�Ib�
����/�xlr�x�8�ܜ���nĲ]V7R��B��o�R����m=H�����h?�z�ŝ�5�s�5��9�^x��I)|�y,KL��Z��R;*���WPr�1�^����b)������NĘi���Ӫtiâ�@<��;��F?N�К]qT���(�6n���~`��`���Ak (~�N	�1�I��dOך��(z��U���p��ǹ9�A�m�ʴ�37+4�.�*��d}��T���Gy���-!O���P�(��r��XZ��$�t�Ŕ��z7q����~߬u5����HU����'�<��x��Ŷ�<�##y����\�t*�e�Ԏ���s���Q��O��w��J��^|M|��A7D(��"�I�q��-����64�Wb��̥�}(H�v��|L�t��p~$�ڸ[���oՄ|3.1��0��풘%��S��fK��GW�ȡ�*��>(���l�</�JS\o�9�V�۪�񣫩�oָ���3�3���Ryd3��
-O��o
fKA��y%��G����@�
Q��Y%	}�_�i�v^��V&��Q�|�K�&-7_��n����l�9�ڹ�=(�qn��7Ux}�)��7�S��Ȁ8��Ȳ��vEXS�d��zJ�+u����L۳*����@`�O6@��g�e�I&�PyIg9�O��q���rFv� �6t�	�~����N������yv"'����$���)�v�,jĳ�gM���4��TkT���)���m�s��4-~M(B�X�j�����
H���t4�,2���NH_��=b¡�N�����e=��4X&q6S[
�X���)M����?�!&F�ds���=�w�P�EcL['�V�wb?B�v�BFI�a���>:!�q��������T�Y��smj*PX£0�t��5%?��I��VD��g�D_B�\U6k.	���Qq����Z��f�ۥ����p�����yb���X��ʂ�+!'�Qm�ށ#��|k&�׬f֝��fk˫ ��p%z\��|�}Z?Oм��c����w�7����c
_�1�ޞ���ܓ����0k��aP��$֚�ȅt�Ch�OB#[��8(��^����V�Vž�]7�ҐT���`����鳞�r��X(�Y�f��k|YB��*;(�(�m���+J���v��	��_���g� �gц�����u