XlxV64EB    29e4     c10�;&�ʿp.W{R%�l�� �u��jX�}�|S�YT��;�л)2py�5"GQK7��J"��:��s�J�#�U�?f&�Øe����爻�0��l=���^�J�ӹ'
��>�x�"o�ǂ���PN��H�X ަ1�"i�'� �.�Cq��,5%�N�a%J�b���Q��s��鰓;�h���jh�U5$ ��'�o�R%-(�ԭ�r���D�����z~U��:���]^z<e*��;+U���J�i�f����ۯ�	-�D�'���������I��.��qa��wd�h�������+4SX(����/�f��'LB�z�� ���,,�ki22� �,l����p��վ�i^��z ��G44خ\��C���Gmj��?B쩖���y̽�ꪩ��>L%����c8��TlT��L��_>�ϟ����e���&DuB��
��0qUz��z�  1t��<zD�8�;�/E��]W1®�B�-%;�@�{v4	�`� F��!Y;l�#�o�QGŤ_�W���Ě-�vWXmi�W�ܣ���)l熲i%�� x��;�-PsW��s�2��wt$����ͯ���⮾��)>X�#�}�)bs��/��	���߱c�\�8�T�=@r�f[5�~�����'�`�����ʇ�%
F(-�8@�Fm�ϝ5Z{���ː1��(���(V�˺���'u˄
�X0�x)�[,�@��8�&8�~��{P4�2͆�i�F�Zb��n�߭�[�nj��!ϝ����	�5#D�Xs�n�8y;x�]�C����lI���C�܏!$�f8��lʤ�p���Y(��� �����g�t��7Da-?���|o�������r%�}O[@�Ն�\*˟is�oU�A'Z_mG� ߑ��NMJ��ER�Gu�XO��!g��!"��P�次z��JQb��8"
t�[V���n��[W?\�N�a,�:�<����T���S�,��u&���m�9$�g�s6��F*�Pɨ�g���N��4ϕ�n!��,�0x4�,���0T���ɻ
�t�%ی��b�>8��t�Zg[;�n(J��vC8��2@��cr����N�� �����[k�&��Lш����ِ@S_��2���g�8���[� �	l	z�0�����H�Kw�n�;�y���Y���@�z���fS4���1�@X�g�ע���-*���
��������;�fr,䝉C1��Fx ���j�%�;��Y���}!={o!n��w3��F��R<�����W	��&3��&��1VѼm0��t���mQ%��|ٱS��n�>���=$F
o[��e���;�����I������,5v;�$"���0�.q�<<ǦK�}���Jνs����^`���#uh+Ԛ�o��F�ns1��;LF� 1�X�l��o�닾T@�û�g= �S��˭/��)��eGȕH���}�I2FQ%�3�s&�i�� �"ڌ4I�\�*��P#`���׍�p��H�n va`KY�r#�j�)4u3�i9o�u��rW{�A�6�j!�u��מ���ӱ��s�-5�N9Υ�^���E2���.�U�g������
�����7Ǔ)��6�S�$���:�AD�o}�]��Z�x2�d�����[u��qN���*��	�fV��*�*M����v�=|\#��(i�^Ne��<�OB@��[����Ul��l��॰��O�S��2Ĕު���Ɣ���.�]x��2����7/���1 SO� �7q��{���+T��:}��fiT�m��G#�G	��^�tdm|��(�^�t/��Qt&q����5Π������?[��*��e
���Ƣ��6YW�$���g;\W�yI[}^&��c{���f�`D6Jz���#��B��~cTLd^�ؓ��Q���H���s�Plch{73�Á ���yZMm^]4��p�-�O���aQ�g��o3߳\<z3&L���Ũ�$�4�L�����*�ŭ��6 �����al���u*�σ�b�IHBC���o��ꊊc�L�%��JT�xD�����$MkA�Pw:�H7��f(���� 7�*���4%L`�D�h�\
�cL���2��wǇR�#A!�YN�<�sj��s�f�I|��n���d��[�/�p_�
�
Q��1�%�BU���oAu�-���>�@Y'NS���!����<ǎq���= =�[�'�j*�	�Fa�[?C��%��ի'ۅl(��/$�v=�峳c��c����/�g<?���ʙ��=/��w��ŜQ�;]o;�z� �E��fH�#�i���uK����y��/�C��y*ؖ-��*y R����T��@��1��ZIzU�Ցsٿ�}��	:�Y���&�������N_[HSp.����e�ք�hd����\t�M���+y����dY��isW=�c��P�'�����6�9�z�k�u��7���|_��!�4�`�j��,�Ͻ����6<�D)#@��ug�y\����4��?/,�3E��Dp6[3&Õ�b��H7A#�����YMl1u�u�� �����$�������8�퀸L`���������g�~�ٮ�J�g2�-4Į6�Pc�CfV�����pPI�V��o�����4�s���e���Xɶ��|���2�y b���[��#���u�o0#Z^ڊ{)3��%_+��WD�ƹ�~�9c���M��Y��JLw��#���Z�IY��́;Dp/ø��䨺�w&�h�5�䨐�7�� 7�������&I�0ģ�E0�\�5*�C��p�9�|xc�p���}���o��A�~����6�_�=��ٸ"'�͚*!��LЧ�}\���ge\���PD��#rv^�]s"�q@t����Tw�>�O���
�pz�7)P�gP�v��-0%Z�;s�Kݼ��h35�N#� a=TA~Gś�"Ogb+�"��T��+#M{oy!��	���%�@r?����h�"`���
ǕT�oDsQЛ