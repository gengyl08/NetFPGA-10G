XlxV64EB    fa00    2dc0B
^����tS�n�t��뭰�Y��!�S�H_BA\�!i�g��R��3�ǫa�#;7Qy7R�	������D�e�ß Մ����P`~�1��'���H��$:��wU�|+�xX5�=�R}�2(�Kh���(��0vG"T���=BD��pR�[=�'V)*�n�R��Q|�Mr&h5�p�%ˈtܦI�H���ss]�������_�kov}�p;إx��J�������Ůz?X��\�Od]�i���)U�Z3� bµE;�~�n�6�j�$��we�EhmU�Stf=����9�($�d.?g���c�{��=S�W��ᮧ5+�1D�<��֎vҍ����'���������+@;����E����,?h��C�;.�N>l�#
�`� ґ��%x��kT|c�(��%��c(�'���>���{�ꚛ9*b`�!��xL��۩v�Iwp�s=q&L��M����PҢ#Y&m�, j�_�����'�e��?*[�'%�����޵��0�2� �-�|3Dr�!9�07��̍�Q#����.���Lm��f�����/����66;���e���s�7�)�#�C�Ľ��y7$�J��IK=�s��h�tq�1��8����u,��N,c�A�h����ˡ-T�m[��5�����E"�cX�f�[�%9?{�6/�
��(����f7Z�<�1*t�4٧A�-��ģ����!/���WKځr��v�æW8�ܘN^7W8T�;ei�H/,W#( 7�E=�vt�P`/��Fm�u�3A9OI�T�ySu~R!�M�j�������T�O�V��!;_2� @��"��G�A��+fP���E�f���au�?L�@]�A8*v�2�E�����e�mQ K�Y<FAA�枮w��b�͌����f'O��2?�_���0}�����y����ٕ#�p����q������lm:�O��Ǿ�D�a��w�!�Zs���rSuQ���K��}����h�ll��I>z�N�/Lk4��=�8�Hb��L"b��U��缎Q�V�ePV(�׀��Ԓ��j�=�0����~�nƮ"��:M���;�1Oo|����俺] �r��+�!��i*=L��O��~4���{��ˈfkXB}ˌ�� J"���sj�I4��⥛�`y��n�!�����1��E>ų��5;Y@z�x��:!�ɂ�#�,��8TCڳVI�H`�zke f�}���`�h߅��G�/F5�n��5������Й��NVE1+q�����7����qS�����i�������ǖ�9KUJ�I�64�˛ǥ=#�i���uĖ��C���)��72�>%W(�ٌ%s�e؉@�vb� D\e�s�_T�Ձ�K��_8������EpA��O2�a�Y�L}��H��K��8Ww?G���n���|)2�3������7� �&W�dK��%�T���q���a4�clVM?ߛLIT����RV�t�]g��r��gG)�D'�T�%���W
qߵ���,���
�{L7�Q)�H0>N*��fz*��������Z��uh��L�ߨE!Q&G����M R��'�i�H�m�S�S�kj�^�]psE���	!��Di�@��&(g�Z����6�~�������]�/���L=�f�k���3��L�ݟ�g�:Q(n>q)���j�{��!�~F�B�����p�2P�HӋ�;�[sJ$���ڡB�2����~RY�_�ZTG��j4l�������L�j�֊k��>����"ູ'�s+�>��efe��<�o"��Lw~���3�F@�'���W�Z�Ǖ>p��{��~���XP����a��+v�.�U
������y�j�	Ʈ+� �Cm~�bKM��;����� �л��&��o2��i[�ּ�&ۘ�� �� 4��!��̌��v����EXG5�Y	M�TMk�ܰ�f��߳�+S���+�<)](�'��֖{F �?:��>��M_�:ޗ�
Z���^������z�z�|#aK�����^W��%���{7IxE1�V����c,�Wj ���{��"%����i��;ː���0s����m }40uTj�0Z1{q�}�7�kb�T�+�� �JF�\M�uq�V|0��b3����YIS�Z�
]٩�l\�k�Q����Sq�F�/o�zd|�Q\�N��	�;�Ȧ�T��N$p ˞�8r���!q����X�)�x��N�8�|)y�8_�2$���+�6�W��:�u���{n8aA��@�<����cĖ�;��]?6�~�M��_�ŗ�t�N�LLqh�M���)�uלf,����`8Ǖ^����>�u^;ʲ�X�>W]����;�����d�q�;�$]� a�w�!H���U�~��[��mn3�?S"m֠o�Mxf�P'YK�ݰ���^��D;}٥l��m�ڏ�rc7�k�#�A��u�:�E���*���� �<go��U�V���B�AYY�dJ�Asքh�B��-����Neѷ��w�0��#t���g��wS8��D�@K��)*<���г1��`S��ϱEV|�$��_kK��;j4�=S^*��|0�n�ѵa2VF#p/M�����o�1�Ma��І��jT'�i��K/B�M,���P3�/zV&���N�!/��"��<-/Hs����:ȡ�j�ǙX_@�跇�N�D�e�֏*��3��1E����������x�W�|�5����尖�8(ީ;�7�{�s�f��b4��m�Iv�`A1D��T1�U��
-~:�A�{�~A�q�o��c�q���l[tNP�-ӞXc��uiɬ��U�P���A����Q��m��*+���3�<�u4I(�Rlcvj�>��4,~�b gXRC*`��N���<]d�N�r޿���	�//�]p7��ٔ)8���F��t1 ��9���"u����!�Hd[� ۹����]��X�~���S\�T~��Z7�3�+��[!an�|Mͩ���)��=�p?z�0���g!4cp��H/���-u��o3�Uu8������&�X�p��	k�S���4���Lw
~�	SS��㾩@lȭ�ϡ�������"W��j�E*r�s�-��[�3�Ic��@zx]�Z����y�V�X�[��U�"9y�'(8��*�C�֯�Z����[{��/�0AJ��@���T�⡉�q�e5�+QatO�-�}�-�/d���� ��G\�G���{m�XҮ��;Ș�cNP+E�5�P6�������3E�n�]�����]���	JV�A�Т�J�\�АV���޻�MM�҉�~�O������
 �ړW�]�:&y%�<D �a�8%3 ��j�^���Ԃ0�2��B�K���	�W�`�G��uJdCJV�)"�=����-���eE���%�6�O��@�?g2�A3qe�_*���
�QP��Ƃ�4�y�E��7ĻI�,L�&jۙ���M9�"�wP�~��|Qi�0t�NMӍO(]\
t�G�����傇�iPJԄC�zo�>��^���vܗa~$]�sP��yg�Qj���q���h ����ϥ��jLT:��	�|��=�_w1BS����^�][z����ER�r(�&���AۓBt�,RM�(�ZQ��Y�+i�g�
t��26���^Equ|��UZ��w��Q�q�xtX�l��9c�mn4rJ0�<��t���e'M��@_��Ժ�̦m��/n�=uoz��/sF�r�a}̎�֪�.GzI3%�Dr{j��W{�5��?�@��՘vH��K7��ǫr�ͨw�+����U題VC���{���`0&���GA����W]k���p�m�?�9�ϟ�����s&�����4�l1�=8�r��?>2����]�Eb4{-���*����O�����\�~ꧤAA�&��ü�'r���چ�OX7��ѷ��� ����Pr�!�ru�W�ȅx�n�5z@4�O��-F6n��6��*�l�/v�ԊoG�=wp#��k@>��x5. ~ޏޘ
���V)�d%TvJ�GT����_	��n�+_RꤦEMq�_��-ʣ\"^�����$�\�IА���k�8��oJ�*���4�a
��&���8�{�Jk@���T]0K	�3�d�-�����RL�ٮ�Sj����[T���v��7}&('|Z婟*\bs�@)��e&dq+f��
�ޛ�(��M�M��j���\��x�ņDK
��2X��ߧi��*Ы�h�����_�9����1'/�M�!�bv�\l�~�t� �"~�K�l�oIT����~��M�$E�W�}�<6?�����,Qd��%���`T�:�Y�mrW�糽h�/�dN'<r����� ��?ۿ�����,>�CDr�����CBr�4��tY�~Ė`⎠C��&���.H�rt�&�
�|jvo�L��j-5ǖ/o��н�1��u�U��@�d1ج���/+H:.�LϘI�j:9wi���y�i\Y���C8�bU�?����L]��f�J4�G)-����KFٯH��T�6���*�(w��[ߟ7r���+7�q{m67hLy�g�/�s�O,�zE^w�7!��f#O�Ձv�t��T?-c"&�!��!�5���?���r/�<"P���Ӎ�Y�8�P_3<���΁B�m��`��o9� ��YB��s~!���+5��I(�U�����:�X��*����ARCF�����Mr�\�� 5��G�Cv���ꠕp��O��O�^�_��J��Jb:�������O1�װ���f���D������7��9�w9�=;�cI��N�pZw��!O���[JF|���\i)'�r�Ig5�.9��?�
��g"�z�&��ͫ&�?� hF�\�XC`���I�`>����������'4���:��eW���p����_^;�2۟��r�o��}�H3��)����h���yE����ܑ��<��HL�C���Bd�{��u���y�͖V"��Q��)�TT}'�.v���p���,4ZV��Y`�w��Ո��O��-06�_J�@��`_�I<)h���#��#�U�Q�-/���"F����m;yu�G"������?�&̟N�{t�I���o�V�+��h㓂7FzfL��m�#;�<r�V$���-�m�D��O������oR�y��<�i�a�ڕn��ޣ�d�X��$�����A͹�y�(���R������9�N�!xV���q���C�*�"���0)��
#o�7��M�&�-Ii������ҠI���I�7���#e�vm��S �r���B�0r��f�d$/�B�A5���^�ᰂ�M��r��JA������/�<(�]n�~��JQ�VF��@�)�ڝ��C���tQ�bPQܐkaP�jr�%Մa���{�|�K�#��@��r|y��	�9l/�3m�_���z]�ǖ��m>VA��?&���K{�ٟ-JTy7Ý��=���S�'�6��b.A�!�&W��=�pOE�2�~d�|�-2��}p�ҿ����ץ����́��;az�Y��V܆$*ؤ�J�� �h��W�- ��k�*�M��ll<�%a�a.Yb��nm�+�B���ظ~P@"{˷�>�q����\��eX̋i�>@��}�ӏmr4u�&���+D�������Y�A����!�?ޑ���t$EK�n�)��<�P��hj�7cWн#�lBdQ=�/j�T@Xcg.����X0ِ� ��>�ش�7�ڒ�3�I΍<W�u����I�d0�^N������O�Z}�v,X��@K��`>2��ctZ��>q�Y��;9��vy�9�-�B
]��7������Xo����*쇻"�;(M�dM���l�yR�+�4��L����dR���f�
.������-L_��QG壋�,I��l^�f��L�c�"lC����_"/Js�	��_9�
!�~P7X��uT퍀�񔕘f=�;�f�.���Oiڪ5���KBa���.�IT�����H��1:~���Z��ax���P���u?T�'"�8v��<u��XQ��7�����z�u��'v <���� &�&Q?:��5t�wCG����Ư�Qm��f�=���V_��[�-'�m�����X��rD)��~�
��◮�W:��$�+���ja�G�X���twWZ9�kfEC��Ӆ��E&�Y�ɿ?	���Ȟ��©��A�e�۳sp��J^��ś���V�4��l �
~�k?Z �ڷJ/X=����0j�Z�����s��	P�gy#���|ڙ1N��lSC9��g�L�ӳ̇�MJ�V������
��e�AKzPNB�Vy��/o��=����0SHf��gn 	&{M0od-��1��Q��_|na�(L��eדc�"/�A
橘�6�v��W���F�'��Ӽ��/ [䰅���-����/z��F;�і_W��u�e%k'~~�k����>�U���)���I�%��$˫y��_[���OR�r�(W����%*�D�)g�t�lkl�+/`�_�QeeJdt����4��{ur�����SW�;�����zeU�q�&Dj���J�yGaKS��`ۦ ��CH�� ����,�)��L���{T�u�5C:(�H��uޭ��5'h)���(:Gc�����lؗ���=a����#�\u�v��T���'����M�ҋ�Z ܴ����	��L=.���Q
k�qӸ����?د�=��}y�g7͎ۦڄ0���z��1���������,��Q\�����Z��ۨ��r����V*K�I��N8�G��"auM�FIP<	{Ĩ��z�]16�A/{z_'{'��N�)�T�f�E�=�������Mo,�T�S$������{���h�R>��/�89�'�B2���j_d[B֫���3Z��<�TS7���&a3r;<���;R[��#ڼ�f��h^�g�B��7���c�9�Ć�<��,���)}�RY��k�$�k���(V�ze��ܵj�����$Ϻ�:R���<�d�(�؂�����f�	 �L	��B����M�V�"�'IQs�-=L
⢃6�VO���Ȯ�l�2�N�0�H��$h�s���&����V�����.U�mi��J'�6��#��#~�d�o�����G�AEq"���7����g;����V��ذN\ݸ%w����s4[��L_�o�K�rN.�:e�������p:���Vj²�gֿR��gQ(�Ő$^2e�ods��Z(���op���`�qg�P{yZø��GՇE0h���H�a^/��e��xb̳���7�SH�$�X�Dwk!:�5��길,�@AP�X��to\��x@�Ī���<z�kU�[��2��V����8.���1�0��r_�Ye����L��5aɱdf��r(���Qy��4&Q�m�U�P�?I�06�oN�B�����y���M͵{4�ԙn�ff+�����<�1��x�n˪�mGuX�^z��_�!�����)k�8&�H�O���)�w�5C�uz���&j����娸 ��$�d������<�&�z��_���W�Y�œ�Ҧ	�'u�����y܋Ǐ���ev�zl��E�����#�����Wm�)~�h�uà>8l�q�ߚ�]����c�_g����1�:&`��߬z^�t.&y78v���9Ս��1W����G]yNff=@w$h�O̼T�����@��rN�� 7N��B4�A7��Ub��4��~h�h:���w(9k�%I���l*^'��g�k����t���s�I�NP��ة b���~���9��ђ["\�2.X]�;E�'���/K��ڏ�V,���dV��1�� ����7c�>���m nb���_�\�G;��9A��2l��\� [sL�;�A�n�[��@��-�"��\�D�Q�D��z%`R��3�V�A�4�6!�����*�����Ӱ����e�M��:�/�~.:���`��hVc���cB�$�@,���]=�f_�T(|��ӿ%��`�uy�t`3g{37MT���*dƾw�3�@F�sS
%��S ͙j���ٯ�e�oT�`�5pTA��q���#$�'��Bco4a��i�l��I�{,���T�D�ݓ^�@@q	7�Mq�	�Wm��]���f��
�%����OGY0�e�K���~���g�����l�F�Hc\���Pє�?z@\�|v2����������T6)o��;�Z�x�����`d�7���/��|��f��$�*'<�N�\+.Vc��_N��Ҕ<8pg��ctqUmD������*�xE	�P~J`S�$����G®�Y���������m�Y&�
�P�h�~B���2eJ`��ܹ���;w�J�-����~F)����o����>@^�Eeߓ?Dv���u�B��}9;~�'B9�H�Z��jT��%>j�a��?���R(�q�I���-���ʻ���d���w|`�O�\P�wmh�k'n1�1efG5�UQ��l�18c��`�NbV���d�4�(]�7שmo�5�NoL���qpnm���"���b�J\7�J^b���s8�`C���7;l�|�΄'	mF0e��Hc��s�/g��s��!�l:'n�)��ƾ ۘ3���N��'f����;�Z1�_aVm��/�}n�&yI*�K�V��є;F��i#4w�o?:&$���TŠs���*a[�
�8h'���V�����#�����YR9�E޸�I)c����5�ʘĝ��w�I��D�(��"�}��q鼹Q�rU�G����O_ꉭ����@���%M�KĢ��g>���<>*��rM#v{�>�Zǻoȓ�+O�)7�Ku�J�9��v����5+��i]�I�8�p+����J˕�1�-z��9
tUt%o�NM�_��L��43����	�)�ѧ<�<��j����*ԛc�H�+�,�����^���?Wf�����fn(L�Ǔ�"�`�U�3b�A�x@�9Ⱥ߁�`�sS�="�(�f���'�d�tx��R�f����b�Ҿ>�s�z7ф��K1�|���6�ȓ��QM@����;��uuJ�
)^>qڹ��#��8x~�/4/T�,4������x�d2����̺uz� �<�]F�<��h����;%����b�v��L|��V)�)��D1��O�l5��ԐP.5���R�5��ʵS_p��b�b��/3�D�\���nyTG)Kx�O�5$�������T6A��}�L��Y�p�1nB�9>�D>9z��**��1ڝE�o�rpl��~|���|Z'�,�S�A�<�-ղg���d�B�x��&�3x�<�7��
t�i,��Z[I�+���u[u�Ђ)�,�$`	Yj4O�o�O/��p�$���"~Xm�vn�=<�G��*��?��8�"��|ƌ��>xܣbyk#"R�n�)Mp�z�(�q^���/��������.EqV�b��
�ǫ��r�M��, ���N6Ԫ*�Hb��t�6c��57r)ej�FP4$�GV��y�;�Nw0�?������W�놑�@n�e�B�7�[�s�ڔz�o��! ��4jb��T�nŪ�~8��h�d�&��졞u�7=��~��Z�Fk���p}n4�#D�Q�L0�2� �G	�X8��]�A��ʰ��z�kS��G�@��W,����bN��tu�ahxN�-���]]n<�8�]�CQ���p���٠O�+��i�QɣRd��o�^x����߀m@2�Y?H��v�]��������b�2<a@eM�?�K��`x�cg�\5*� 5��(7���P�I��ę��.�� ��؟�4a$:�t�]�8��� 	,�W��11(I�K[��k�E�X�?�^�'fб�{u�+����,�"�0dR��H�6%mP
,��{}|1�tL�|�ɢ2脿�~݇�w��h��<R�Jf���x��h��351�9��1��~|����h$
�W���A���:�����jY*Y+�ٰ���=�N�6=��Jzs��T.7ao����RX�8S��<��:�r��$F�F�a�F��؋[$G���aϭm�B�⓴;v�Re�������>�Mɥj��[�(`��p\�&��L��`U���_��(��ƚ`>��l'�����mN�D� ��N���Il
����3�r>�N�؜o���a$A��FAǩ�R�L��>��ڻ�mJ�VI�Z/����{R�"k�3��:�J����X**~�2�=�Z�X&��CCU)*.,�����6�*g4�B����x�Q�m��<���j	�?�B�̠��4�坰6�9��Gң��z����NB{fU���3������|�m��Pq��*��$���Ş��#����� L���{s�\��l��m5-��梄.����m֨{+�b��Hl�/˿q��*#��a��k����7��x�R�<�%���P�^���TL>9�[
��C;`]GH˩xZ��-��s���Y�i�,�Z�7l�a�r3�<�M�Xt�����Ah
��󡎠��z�ׂ������#�.@��gY��H�4y$��W
.�y6�"ãp�
��5Yfi=iOC�0#�+ܚQ_qg�Ҋ���}��n2��G8k��D3��A�^��nh����
6�l�����Z���1��%,��a\�N�cYV���G2gЍ�����Jn��G�=+�@l��d%ᅐ��f���YmIM�<�9�𓂃Q�a(5 1����[�@-���2M��c�}�Qyc׸����́|� m�}�Q�c{��T�D�*�9��p�h��e�>%f��.G1u��M� /'@�/�f��
��HV���4�"�|�����bi�	�Ix�	���:ӕ�"y� ��d<��*����q��j9��Fo���D�o3
y{�*�Y˜[1d�	ӹ��7����6^W�T�Q6��'G��S#���dI�h�ޤ/,Y�d^= ��z��mzg\�4��i��H�XOO��N���鮇�>�/��؏$�;Gz*����)�3w�f�Qxn�r��}�NсP�
�bb�ҢH�s�Μv��ȇ�]��'`	���e��K)	2�ι?1�9�j�a����h~L9%L�qx]w���Zs�kA��kI$���hȝ����ʜ�2>��x��XB3�<�R�+Y?GO`]՚�n3`�b��O���-M�-(�|���!���p(&�������lF^0'���������W% ��Ae�$v���Ш�!&n��v�G��������V�&U�+����=��C�a�fo�.^�*�!v����L,��*�/#�V�	�g<��ٖ�H]%}�[�ն�T����jH9Z��h2�M:JͲQ�sQ�ʲ��A��qi0�P����oeĭʎ"Y�:}+�O�s�DP�؝lօ���J�^*'ZL��a�q�b
�1De[�"�n��1+*�p��h��}W�Q�XlxV64EB    aff3    1c00<kE�än��҄%�ڏ�b�w:X�Z�� �<���9��}o&��8
��)�Z*-�A�НS���x)̧��_�vx�B��ǝ�k�V5M}U�Ι;���B�\MHE0�l*"[ɩX��k��˴�����Q(�a�kN.�n��)AF���Z�� 7��s���/�u*Q.Ψ�����LC��i4��O�뱚,��e�ʨ:*&�J���'���A�~����7�#@XS��H>�������71xe@�X��xM��3�
O>+1�Я�(���0�Q�	k�P��i�9���\Ղ?��m��Y���?�'�����ɛQU��ٿ��\Z%1���l���bj��j$�O{�!���K˙�.���2ݹ$�_wM,p7/���� W&w�J�����K����Iy�Jv,���qB/J�7t��2�x�h���:�W��M\Dc�&R^�1��|~����3�8�u��dP��e��J���|FlP��$^�>�mz�GN9Gn��f��� ļ
�{��f�<ծ�Oi�B��G�q5��̉Q`hB��|�+�Tz��VB �Ǌ櫮�k/�a�����哫
\��5(�'�q�^�2C��f��{I�M��<J������?qnH��@��ژ������qj ����.O���:��!n�i݈_~�/K�Ŝ�z7Qj �&�\xg3�� vPh���L�F����e;�{ǦFp�s�sM��F*[����5Z����\�>��vH耤"��2'c"9K�c�I�r���;��OC��NSNPP��F���������y�0���/��7�6� ���ξ��4	�(�౏DX��e���#	�i2��i�.e�%l 1�T�L-H|I����o�ԯ���t7UT0���������"�3F�R����`�h]G���Q���Z��|��{�`����m{E?�6�����T��{䕭o;pEM��o���|C������P�:��-�T�j#�q�۴D�Rb�Y�qYYc	�V��J��0�C�̴%o��X�l�(�5��'��qA-_�Xp@��6p����ަmH#���;�#b.P��?���HL~�@��"�2��?�F�`�5���֏��)dN=y��/���U<��8��db'��g��[L�H�|��1�V�����]@��`��w���S�\8��Q���,�?D�&� ��E���T����+�i��w���a���G�\�k�ԽA���Y�\��y�5��%@C���8j=p$��ۉ��jļ+��3cؤ�����S��I���dF�p�6x$�c`M��ᘙ�N�\oF��j�0��.C3,G�[��pޒj���.��$�"��[?ဢk�by���2���ҕ�e!��<ƥ6wb��l'�ʰ�K�������K4n�Q8 �W�q���SLk0��f#;�:�!��{��M���+��v��Ad�僮hߡT��j�F��O��T@�i�6>�&��-J��'��qDj�a�.˯9�
�6%���ehBcB�E]G����_�����b����0��" �6̯����*w���ys�^�a���_�-�h�;����m�g�[B�a����С9���_���=1�{%��ﻂ�_$��N�ⲡMY���d߽wF�y�3�cSs)��W��"�,�m}�0�X�l�7�K�ȯ�7m$M�!���8K�U����T�g-�
+����LJ�G(��r���g���5 fA�-D���R�Z@�B��$]<���Ρ?�y��OV/9/�w����c��x=r�z,�5ց�~s��f˺a$��Ө��B�WN���b6�z)1�f5���q�7�N(�8؋��Ƒ�7��o�-٤��a��͖q�s��-��^Z�>9�7��^2�����;V;��	��w�B4@:�`k�^��n�{4
��{�<�1��t@3;̴`�b2&���P�B�eS�Og�$���9�:�M�S��Q�#�Þ�����mooF���
[������P^����D�G� �����G���ʸ*9{�}A�9ko�����M���A4�J�Q�!Ӷۙxۀ��ɍD�͊ ��7��Yx?�2�u�ţQ���ȱ�Rc�DG�s��ۡ`/���4��Y��n�V�ͬxX�.��jy+`US+���!0���E�\W�g�uL��0Ll���Жp,���gi���M��4i
)���5k��}���P��*C"5��W_kG� ӡ�WF�z3p��w>撅.����|Z�ӹ�G�>���O�L���5����~#*8���Ǒh�+l9���Y�<n
��.�6c��O���+����!�Z�ǽjM�� �2�?��qC(p9���sU�a�k1f�U�mP����-!K�b-:I?X��尞:K�Rl��bC��mG�-He�j>��F�G�c;�֦�:T���P��>���<���Թ�zY�w9��>)��4#��V7e���/J���3�d�#(������z��&l��R}� <Q�\�K.[�'ۚ.J��E��&	�_�]��\�.ubƦ#�6�r܆�G]t�����g��%Rk~��ea�k���_�K�:�i̻i����������S���
�&|y��p��q��_��ן!�0�������_B�	��A�Fu�8���]�p����@'��D�9��6�7��$����)T�v���?A�n{�yѵ��̱Hi�>�h;����%�9��?X����k�@B�33��#�Rr�((�L+k�j�nHL���j�K�$^�S��e>��7���Ӝ�/L�4_Cb�}�r�,�p��!�/Mi����0ں1�F��\>�?ЮG�,�H���s��M�k/��t3��\��7��=E��ҥK�t� )YH���������GQ
�w-�8��RN �='NA<9�Պw%�B���|k�6M�Q����9�k+ ���e��ͪZ/��j%�Pʧ��bN��|ָʶʳ�kv̈́]u=�FXV���LJ�8�&�ԉ�)��x��#9�q�t  Ş�c�+����{`O�����7����g��|�Z`�sX[�(z����{*G]ǻ$0R4S�b2��b��c&���v�cvZ�����Y����W��QΥ��z=����U]/��S���-�)S����Z{9ds4�-KT[��Ar�S@������������!V�����8ӈ���R��e͵PVC]	m��9ǵ{1��0���ní�C� �Ġͼ1���'Ɩv
�vohWO2��MԆ��`T����j�5#��.��k��,ׂ�疮������Sm��a[c��_�)�O����_�r��L<Qe~�>]!ר酾�p�}��s71����d|�:G�%��X+w��?�lN���y���D�򕌬���Z��|+� ���=0�b�����9բ%Y�"���v��,�W�Nd: �,��a�mT�D�/��n;��RB;���Af���+6��s���Y����D��ަ�q�.Q}x��؁��m��69e=�ځ��!�{��鷣�bǊ�E-�	��Wh`\�m[ۛ��R
M������=��Gm�Q�7ȫ���
�Ψ�芁`@���g��R��^��S�����l{>G���V�|3���Jw:�����THA���R8��8X9\����)��m��!�/�
5�#plwg:�-#=7�p���x-Tl ��]���IWH5=�o�R�EQ�N�Bb-!.�@]L�i�l�dU��|B��4up8����Ȍ[�x�wd��QY��?�TW���&�.��W��rυ�%��f7��X����$�@������C)�p���cd�/1
R`GS��*�o��*�Xm����ʏ������T5X{٫~�l�F\�ik��ײ~a�)��A|�!�^|��q�
KL�JO�6���l% hxM�Z�O�.i�]c�Ei��#
�6Î)�V-[4Z�cM��^��*����57����!b�(�3e`��󼊕�Yk8�GP�����Q�H�=��"[���D���^I	�s��?����x䝗���-}xtZt��o�W{N5�9V�55���N����e3�Gc'Х�r��L�"���h�gŦű~�_�'�@�1s����@!/Y�@`8A�C�@����=�RL�e���@z��i�%̇�����,;�@E�' �86��n�<��,�c�	�=�f�v���03���2�T���N���B��w�%}J��)
E0����a�revE�z/�W��{q4Ns{��ʧt�lj`�w�Aς��9	��=p����M�)8y�P0���G���I��!��6�7�(h��]᫨�E�ి����.����p�̈ �=5�E�921��W�܁N_��(R�vd	%�
ɰ�K\K���Bg�8���k�x�Kh ���nK�E�ҵ���}�����g^vok��4���A�)�ql%��t��Chz��j�<,%��oT�6��f����`oֶ>�BL
��Ɏ�d��r���$�����U��r����2�SN +8�
����	�ҭ��0�Mg�, �ɲyhᕢ�����W��	�Ժ<�(2zC��V�<�9�_�����m��?r|H�����YN�<Sj�*=@yO�pޕ��vj[��r���KG�P��!��ra�ڮ2�!�qg����֫Q1�d�X��
�;��K�狮s�`.֣��m�!4� 5�z�j�n���֭s+h�<��W������R���@-�k� L�8�?�5H��rԷ�b"�mB3T7�:��#��S��O��/]L9��hc��m���G��7��g�iw������{�l@���,������3Re�`�}��a���`_/V7¢/[k46G�A�J�,�?i���q�h�˼�i�I�<ܺ��"�T�S���ɂ̲�m�|c�;M���Д<iJ>MIz���.�=Q���&9*��Cq�;L�cz�saa
W�f���>`�)f�-�He�C�þr{��ਖLD�`�P6�4���U�X�����6������O�W�-�'�Bf���hݐ�gb[5ɡ<ZW��FT��݀�cC1n��mc��$�q~���te���r�{F�{���Nb�[�8dV\r{�ɀ�"<��t_�ݏ ),6V���
DV����ᝰl8���P[ �i��,6��H��C>�6S*��gEӴ�F0��	)o��U�b��B	���֜������u�}�@E��K���N�#���G*�T,�h!r,��R�v��YxQ:�?+��$#��nP	K��,�*e�tij��|�"EE����i��ͳs�t����"G�턹��W�_�I<��K���m�1I���ٿ���L^3[�Էs27�d���w��#J���Q��YZb��B<��jvٹ�S��/U#�D#-BRLf���I��b�`8G��*�\f{lZk��~i�YY�0<�VG`,݀�o�v�m��F.��5��͕=V�Y�D�?Hޗ�|�-ᮜ;�y}k�0��-s�D�+0�8EGy(QI�՞W��!j��C�A�Y&����ҭfH1.��П`������B�*��eC�.#�>��������D��?|���k�{����`�̙�XyN��KY1���a`4<x[�"��Թs��҈�.-���k�zk�h�5��%%���2z��.{�����]���h/������wY�m�]?T�S�ߛە���D_8ν	ߢ�������$� Ϯ� �QHN� mɝo��6�9��;���*8.Gn�I�+%�<��o�%�Hx\�P�w�^�~�2�ZH��%i2E/��p��C� ۧ��C�Wn����ᗄ|M�QQ�z3���R��J���:�i�|�����л�lR����s%ƵO̿$�V<R��DO�YV�R�<3�x�U�VE�{�/�#?�W�}Vp�It3��:֣�:�J�Px��
Hw�	j.�����2�P,r\�y-�|��5!��v�B�4���r>Q��Ę��_#0�E�3���(IݤJ�&��Ւ���'_�CŬ�Y��+}Ax�N��r5��(��7���zGǬ�"<[_b*���_�t��]�����K����"�_���Dz�H4Ǵ4�c���6���N��;��-����+C�v Kȸ�e�[��3�5Qp�<��:�_[3�]+�ZF�n��*��"����������~_/� !=������:�4�$l2����O�/�W�P��T3�5QH��Ɏi����8i�����L�d�������W�M�<*��}����OW:.d��� �pcX�͍�o!���>ڪ�����\�,O%�O���(m�{��r)M-�s��Nm)��,��Y
,�S�"Wo{S���5��H�V�MZ]a�������2侢�Vn(�9��^]!R��j���#T�퍞���pۈ2�������%�&(?��[]C���<�q<�Q�ez�yN{�Wčv�/�����6�Y���[�t��b�-
��.Q�DB	Wtˆ?�h�:Ul����pAQ!A��0�<J��
��eY�/V*���� ^hz���!X�-��/�{� h��T�Ǜ��%�g`�)ˆ��%���wMj�Ψx5�O*^����t��Z�&8��=���K�J۩TV���ƙ7B�_��}r���1sJ��/�֤p[��2q�2���?Ѭ�x~�0���z�i�L
X�[�?������$n�5y$������xQ��8 �韡H�mSF�P��OJ���#+�}z�RI�M`����*>ZT��^zb�1�ز��*�G��q^�
������C^�)���F�|��*�Iۮ��U�Ax6gH.�k�
(��G�o��{��$$9T�k�Sm���ډV`��r�7�2)+g��}��f&��~L�͊���q�Q��'�o�5֭��i����[����~�F;H#j�	�d|?�ʫ���w�|b8�+s��W*��L�K��
��P��*�TW��=M�]b,U� .��Kр��tå_�k��?@,м��Ԃ+�w7����I;�Q��Fga�S��5����ӏ>~��b��;�