XlxV64EB    32be     d40�J>��L�Jͽp��Q���H��?��6�W/����yn���D������ ���
VS���0���lM�؉�����<�Q�IϓS���/��:�ᔅ����,z;�׋�N�[z�U��	�@1�xʒ�$؆� ��8k�M٥��H�4�E��V}�	�i�q�FNz��du�H��Ɨ�����OzK�t	B�o��D�������X�+���H�z���䶝צÐx:�-��FX�x�)�o'>L���4yt�~ʺ�mxK�Q%&�囄o�Z�o��m�N������a)�p����9�g��p����5����_O/s?x6r��m�9:�5�EM�v�������^9���h���0����wh��cw��P��a6b$a ��3ȣ�?�(3^���p\�nq�a��n�V=k��Q��m;m� ����m�Z6�f�R5�,�*����c�f���	�%�T�?�Y)���A5�T�Y�o{K��&0����@cm�^����z�l��G؜4=h[­�6V$=�8�,]Y��r�j1�K�L���6񴈗��`����qL�E?���E���B���ܫH�c	L������[b�a֤5�Eü�|E�p�U��[wH6N�%qj�H��ǚMU������.3O��G1l��@��ࡖ�K��D�J4?��<R?K� Ƹ� [?����_"�`M� �+?zZ�v81���$�ݿ��R5�V����B���kԖ�¢�Q��~��2�6]���b��� v�K��P��n�9�W��R�!�d�'w�2���G�O�O�tE��㐫�,D��i��xr�X�O�D^ﶦ&�4 �X?�nw�LI���g�`��7�z���g[��y��>���|�$���^���0����P*�UпA���wB\X˃�ӓ��"�dQX~�1��OJwd���+��3�E�
S���&��-��{z��6y�)��{�`��a�,�ջ
��e�fZ]tO)�*�����������MH�?N-~nS���/z��mxwpy�ʂI��L*��J�	��P�*<�|o���(������׫3��I�6&����_����;���^Õp��<*��G���pr��W�u3�m0����<%z
g�L�j4���m%f�����F��g�Ī�ׅ���⽿�����9ǌ)�{5���ݻ����m�?��s�l�9ܰ'?cn�1��h���[�	�$S���yz�p62��v
q,��o���'��-�f�3ڱ����{�v�����=��9@��P�@#^�*�h�Ce��Jom�����v���S�w���.��-�f
0���O(41a���^����Ӑ	�W���Ն��?k0$�z
S��ZQZ�ߵ�7�g��Sd��c"�o�~]�P�pJ�?떛���Ʒc�z���8�˖����Y���$A0���1�֘\��6O��{����]�S����㝨p�P�ʹk$�
8��1����z�/>�#�\+��s���\�|}��]ApxR��7��uYr_xTf� 8�ћ��<�|��������UlkI�����]@�����,t����h�v��npe?���.�j�W!C��X�qs�Q��x$'(���CT�!���s��S�z�!�ו-�|z67�'�����y�<sO_�QTr���A�`o&(�ȹ�����O�햭̾o�H�ϧ%{XD���[�C���>��ȱ�_���x��cx�6�f���: C\�곐����@�fw�T���A�"��h0��4�cc��)����l��c�����t^����ge��YR�ӷ�y�>mv ~��D{6}�����;�w������~�0�����,�����'$xi�!�h 7?}|��|߾���}-����i��0;��{�[�E�	W�z�TP���aN�H+�J�"̂e��;_0� >vb��REg��H�?�
��i&�]v��:�VD��Zv����ف�;f�k���{��+u���R-����9򒁌���z>�\�ø��Xk�j�v}�#�[5?��x��' �D]4��0ڌ�]��P�H�e��F�=����^>�ߎ���.�F��zlN=x�(�;��$�?�6!�Pԍ�J��)��u�~XƇ2�#x�;!f���^�Q�;�nT43�f�.��� �|F3�ݡ�*�����eV6
IK�pj�	
s�9^�PՀ�a�ȣ���"�C��P?*l��.�76�7�^�6h �z;[�m�_��괩(�of�b���8�[5~��S&/�������IE�������[���� k����*�b�w�TM)<`j�4�
eKU��Z;O1����/���Lr���ee��2[�U�ߩY�a�vz��@�{X����d����Wa�LO�uDq�����-f���y�p��� f�t��1(O�����(���q�D� �� ����ῦ�*\Q@��V,�;	�{���_G�e�ᢞ�(�v����<�Wl��)��Kf'����t?�E\�UbTav��d��\Uq1m:"�v���9߀�H��"r��w�E6}���\�J��_N���5j�)����#z�� !:�%���u#s|y��Q�De"wd��%^F���w88���4^�ӓf��H��nBB�@��&~� �\��^��g��0:�v���kI���������'`��$�x�ES����	����5�:��J�&�7�iM믧�2���������Z
L �W*��@�)`=�nhvԇ��o�zᶗJ���J��#F�"�m%B(,��,�X9�mJ����}m�hS��wE�ag}���q�s<�cf�gVIi�7�_�w,H�I+n�mW�}�N�ڗ�:�U������W��x�\�7�����jk4l9Nz�k�5�
����ڈ�Wjk�V2=��D�NvέG:f[��]���y�Y�RV4�ʵ����䭡�5�$s����&�G0l�� ��)<6�池�8g�;O n��K}:��VE�����K�q�b�p|�G�3����'��>ηmC�>oh�C�����A�%�@������=����D�*<��lM���6�#ϷSk���;/� �k�lߊm��qtC��P�3��oGs�G�b�vd!�5V6w��w�����6���Æ�ck�۵aː��7����a�T!����I!�a��%cSbgIN�3T�w_]sM�iߺ�Б���^aǼ=r�i�5�:v��K�t��ark�s4?<���
���
���(��S�������=-_�#rB<�xν��(������9