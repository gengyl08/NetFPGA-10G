XlxV64EB    372d     f604�}�8C���:�XG�n�+��^9��\
ev̰-dom�yu=77:�[Ʀ}Чt�Cs3������p� ϲ��d�6K�k���ؒS:p_��B�S�q���c1��8�?!w�|���<	ڦ;+~�]��.1�)�;R�p�J���B{ 	a
��m���0x�¼}�\��xn�o�<�]��nC�����0_��/!�Y^���LP�]�lϔR�j�{�%�|�0�.�^J</m�\6�0�m����C�4��5Hخ�M7q����4C��E�yN/��s�����c��ꑑ��f!0l�O��o�g�Z�kxL3҇K62<��oh� ��/D��M�-��߲�|ќ"s�ؘϐ�K�H \�O����s[Xb�6R����3�����߭����("y�6c���N�a�c�)�Di��=��OHi�D�#�D�M�:�����{�8��x��TE��ڦߵo��������*I�dӰ3�P�@�%���E��a���P"'*�u��V�vT!���>5"�^�Gw�W�
H�jGz�-U�8��+�L~d���F?n��y렻��jF��TE93��@�!=�JPm�Հ6 N^e~>�:uȺ G��T�N���B����Z����SYVZr�,���@�G��Ԏ:6�gO!���b���L� 	ފ�=d���Y.����v��K�&\/2���wʗ�����P���6����vX(�ӡ������[(��\��J�
z����Ce���/H>�T�?�lv���@{��vUѰ@��4��&���WJ�Bn�6��).�q5?�V	9|�0�³]�p����E�n�W?�R���Ǽ�E�H�^����m�9��j/�OfOs-a��O�}(ª8�6^U���ϔU��<7������8��m�M�=� !p��J��{��R����D2%�I,�x�[��_i�;�l�~^4�!���o�����(��kJ+ ��m�z0�]$ ǐ2������W��ڟ_�3P-p���XY?2�3pK6FZZe���V�N���	n��*�INx[$M<��R��@!z;�)��sy[n���D��=R�;��ο�1�;��w���\F
��n�w{�8B�?R��8Ϡ5��p5���bU2V��Ƕ�cp�Q��F6_��'UE�6�Ϻ��ʩ54��m0�l��;�$t�݁�ʒL�܋�f���j"|F9���H��v��V#�=��X�W�h�g~DUA�C�:�ǆns�K��?�󢇍��LK�0}AN�NԹ��<���Wd���UGSc�w���,�7&	����$y��/Q�F��D��>ى����kH
�F��m�pV�e��К�բ��YHp@�YIʴr��f��"#��ת�7����e`��m��6e'��#u�,?Ȳ���֝�eb���XY|���ş�$Rg���1�12�}��2�8�"T� p|X.���W�h��U�G�5]J ���J����]k�p�9>��a�7J�c�����rF�7VV@�ѿ?!�k%y�]���@iF¯1���K�̫z�v,ġ��מY��}�M��8�\0�m^��7�T�#�A��z���u��Kr댡�I�ZÃ�Y��V��V��k�#�<!+��E�{���t����+�p�!J�������� !�̡�ܜ�]h=��F;ug�U����[I&�����j[�XG��F[]�E6PƐ������w�}�&3(0;����'�C|��ˊN��\jnd�n����Y��P��Z69�C�u�ζ�~�m�:��Ӕ܁&��^o��I�}���_�D�B��Ou���ݭ9��i�5���+[s�6�떪�����c>��y�j�֡��Ki��g��	Zb�i���q!�dֳ�.m��S�g6������ӱ/^T�5�J�%��I�0>�����F���������؟�f��<{�ݓi0�T.>�$7���ۣ'I, �ȋB�gխ���‱��n%�r�0]w�wٲ�i1��]����pP���kˌJ�z�H�}�/���o�)m n�u+R��C���?��/��\�ξuغ�%�S�S:�}=������&�D�3�Iز�}��BZ��-�(v]2Ď�i�A���\mdk}��<�D�b\$!4!�x�ƀ��ɰR���w����N����K>y�Y�uֆ�T`0��{6 b�?�c�\�s�d~��R5`�ʸC%�I�x;tZmK �9As\�T�Z�a@���#�Ko���+I^>�Tf���zl��	��@)Þ�8`O7���?ҥ;!:�a��z�?�&)�y�)/�p���Yb 9z�j�̾42��FE׼�F�U	XI�{�~����!9�l�:d�D�m�?/�^�}kV]����e-9@;�{���݇U��p�ng�@�d7��w�!:H?���
ا����,y�� ����pr�)�����ᙯ����u�e5��Y�W����d�##��o+Q�iF��D�
��(��~��f���q] b@��`��'��1ȫN\���F��Q�E:�~�I~����TH�"����C�U����]$�Մ$�
{ĐiN��4O�q�%��� �j'3M���4R���Af�h�q��\ybdf&c��H.^��ψ+8+_�p#
f���އ6 �e�$f�dW����FA�M��X#\6�3g_��j|��7���|�À�2Y��@e�}K��5���%$NQ�i�[F��\7v��j�~�D��\�6,���=���\�a�rC
m��U�������q�Mx|��2����Dɷf�H�1x�dɔj�������K��vD��>8	ba�V�=SA�=�Nճ<�	%fiͦu)$#f����9�����K����N�0@�y��j�gO���j|��Q��H�v; �(�/�t�� 8�����3��X+��-���"��ҡ�����l�f2y��3~	�ّ�������$	I��<��K!W$���a2�ʎg���B��*D�$�Z|bk�z)�3���F%H��cC�G�};#N�MN�ʇ��Z!T�G)���P
��7eǿx�'��'l�)R?�&<��\�ťf�������gq_
"��\+պ���)���4�|k����6c�9`��E�I����Ɠ���E���>[YV�* �ő(WxWP��?�R�M�ko|���{�j~~�]���oܫ���k ��P4�'�R�h�V�/?��(�+�U���1��ݐ������$�c�d�1��JQYk-���w5��A�Q�K��WOG˨�j؊�id6�u<��Q���2�������A�x��'�=���CA�o"�pl}�腌[-s��ؠ��DpKΫWH]k�������o���P�����m|Uy��ѰA�ߑR�8��n�oWƿ��YѺ�ԁ��҆ñA�k�[ȉ-
������f�d"*'�f�� 8Hk�,[�%���ʡ{.��.����P<;"�o�<�n�`��ћ0�"�k�ۧ��� �l�O�+/q��]n�e����)a�%�փ�4HkSœD��褒\j�Z���b^�$��sΗ�˃O��j�Hf*�_y�0K��Ms�����1�Ӭ�Ds޷M6����ۙ�֫)8�A~3p퐂�;�E��zr�a�[;#J��b/t#AS�[��[�y&�x�ƳP����ex9� ��n�7%�f�r�����\!.1��AdJ�ryZlL��)/'h���b�n�q;s�6�.��&���*�NM���Sͩ�h�baɴ���=�jw\MA�qqe�W(�J��8��vTDB���N	�����ϖ0����OvgGNQ�����<���d�Cx�Ya3�r�yÛ�9cx�m�]��+K�6��_�G��0