XlxV64EB    17f2     9a0L�'��u��ki��ǘ!�P�&�c���o�4��63�?V���q��K���f�Z��!w�ү=
�����3�G�`��:۹cry�)~W��-�)]�<��l�.����
x	tÇTa���̣�p�OyЬ�v��Z� �P��>BO'F��.��`ӯ�-c�RƁr%������]V��h<	,�,�gk�Q:ދ�q�h�خ��+n��ｆ�x���0�9���A]I�E%4˰c�RONc3�'��tS3!���ؼ�G�Q�h��B8�䐰b+B�ƿA�,e
�6�?l^��a����⡧)eUQ	H��|��~W�����������!���dt)�i�
�'}x���h��p|����Ȟ����An�^ǰ� pu�/)�����'9�W��	�bN�����y�N�OTnn�W/���A�hw�9��?��PO����_th���l>>�d��'�jicC`��jc)��-�@v������g[��M�5�) w����Y:�,�Xv�R�b�i��T�⎾�4`?��k樂�ꐂ�4���-U�q�v�vq�-[������~<��b�_�m�!�f�{�*އ� O�Q����Yw��υ�붎����w�}��Ӓ�Ҭ�y��D8�	^y�Z  �!1�i��o?��Uq\[����R��w����͗~�q�vm D�&� 8?�+�:[�s���v�݁o{}{���(���R��Oj��Ό.x�OK 4e��[�j�q �C��Q��HQY9Y�J�?Z�1����&����#Z�] 0uG�F�h��Mْ�[���E?03�E53�Ѷ�ؙ�u�p{�-%cg"o���f8;y=�{Z�{ h;�|c|ñ���n��~��=����~�Y�;M��j�)���lB�{���<;T��sY~�uH�4Aݥ�,��V43��t*�u=�f�:��aYd+��}
�\�R<����|�R%AN�xȱ���m�v�����ppU�3�;�"cHR����"+�˓��g��O�^�d2��Cfy$~�)�}?��E��t�8��hP��m��;�|�T���.+���7L�\��Š���e�
`�/�(��u�G�]�����Pj�<>�в��x��&����w��!�7Uu~�{a�o,�ՅK����V.�������U�Eo�����/����\���Q��@V����u�E�Y͇�g�vE����f��������>�'����4s��A{��a.�̴���ء�p��iF�C��S}�U2���ˣ�9�,��0�*����T�Έ�k��a��R�	�Fv'd�/V�w{Qu҉��1��,
v�D��_�3&���3B��6�z˞�5.ǰ V�#����?-�${�I�Sf��;��Q9�gȋMm*
�Tj�j�Hdj�0vq��u�}M-���*�Z&�O�^�L{d�Δ.��S�D^06��o�� ��]�HN���_��|��|���0�"�ѱ�����綑�@�O|�X��b��7��W��0��A����t��ߔ��8��6���0�O��5��݂����ı@�OTx�^^�!�/V��hAK�d�˟e���B�7�^�wVFZ9`�(L�b<�n���q�ֆԀ�v�`v�%QP;�',����߽�;���q%�˼i;���5VB�<���h������4 K��_���U�(ml.^4?s�،PW�h�mX�Ql_c���ݾ�]��j�׶��1׈�&
"j��f��u�Ƽ��!=�x��1�q����ZI-`��x��s��>��ͪ��"�_=����@h��#?�Q~[����e��/�{��P���`�Im�/j�K |�����������Z�dZח�"/b�[rẠ�a��(]k��|�\��2��`��_�7Z���X-	e�)~G�*L3�ͥ^�a�߻I�"�S�D�"���s)f���c�1 |E�Iь���L���)�~"zʝ�,2T�aC�nmK&ڊ��������&𝰇Sg���ױm�$w��B��?�˛��H�L*⊴�j�Tw���6�ܐ����J�1�F�V�m���4������U����M����\a2�!ٕ��j�*\E�E��6��h�$9G��Vv_T7=��0����8{�񘢶�4��,��:��=��ͧx2�8���wK�~��� t;_��<����BHP��B�9��c]�-V�@ yP��j�]_w�p�}��$A�A�:@ �|"	��B� -�O����0�au/��O���O��O��c�Շ!�X�AlP��MV�
s�9 8�ɋ����H�f��?R���u��<v�v:z�s���ރF4�^%7�ܣ��?�Йlv,T �˯UiDũ��]P`��R <8�0�y�`s۔�l�ho�Jk,9"D�%ǒ\^�S�׮*K�_���Y��IW�a1