XlxV64EB    1f60     9d0�rK?���8AM��Yw���B�9j7 ��+��XQ~�}���z��v��@Zq}8�iLM	�:�;�{���{��^-D60�̔;�<.)��=3���J}U*צc3]Kf@�?i�%����%�	�W�������H}W�@������{-H��P6��Iֹ�ԣn#1�-����{v.�i���Yk�~%t��o�n.f���]/v(_2W�[����(iv�~��}<`���B ����J`��#e�Kn�˼��\K�� ��.u;���="�,?�+ZB��K���@�a�H	6>`�|�	��;�d���*�z��QS]A����'	����)��{O�r`�6��W�/:5��K��{�~\������G���Lm�Y5zV����X�ܗ^.�@���߃MX1޵pĔ�1�+F��T�qZ2���3A��yv%?%=�� �~	h�q���>C+a���K��|��4����F�\�$˟�d}�?d�8ke�o8/ǡ���,:�-�"=��Ƚ��_�ߒ:�,�?���b��$9��T��n����1�#E�w&�V�4�YD���N�ƓM��n�ތ�\S4_/�'���/�.ma}��y~����P��gܻu�GC�G��V�1�]W�>�iY;0"���4@�R��k��Y��w�K���7"�d4w%
��MN�����v�P~�3^�����]��s��]�Z�{$��j�K
���F�w�8�F���:FB�j�O�AFj��������sA]�W�m�4�yu� �J���q��֐�Z���e��S�.�zR;�AE*R6O���ABkU����]E�C�f�~"]���aq����P�,t�baq[�������I�Fj-�d����X��y���{�r�.���kq^�
b}A&E���W��:A�����`J�� �X	\�W���X8���us�S�@�rSM�4����D]WEv�]̥N����r3+
s�r�sh���Jm+��.���A_�������>r-��iPGsd�&��6m�Ԏ�dR��8�[H��3A�2�;I��-jj�I�{}�N���FBs@�^	[�>A*��~�\D�x]`hI��i�|����-�j�ʵ��U�z�� ��� ����W5 �KI���GJ6��r�:�Zᚧg���Gd-?�8��^�?y\,��,ԫ9��ve�Y�`��'a��EZ��k,0F& W5���nۼY���yP�nhw�D9����|�����@;e*��u�lFd���/"º�NqN�ރ��ϧ/F��}��2�I�r|��/3J2\Њ~G����醮|I�OuA�8H��aX��G�����\3m�oLNDW��4� w!t�J���^7_G�teP����,޷�z�H���I+�r�i���Xf�`��Z�S7x|���V��T-88x��S�H>���t�b�0�N�k#�ƇP��D+~$?��Y0T��V�|dY�(/��?�t���w�ګ����m�>d��`�KTU�)��>(Z��a�輮�re��\��;K�rBL�"q�`�O����SR�S�Gy��OsP��X6�����u�����k�~OAX���.�-u2�:���jV�x}��RO� ���ԕ���HW��_g����#��OHl�z�(3%@]���ZKtdT�fĿg�S{rR9���v=K{������������-7a����D�{��4��@�J��޼m?��6����p v�9�m;���r[��_�V�}�tx�F�4j ��O�!�AM�ttϞ."�����9=�R�G`{�X���,���F�6(�-��>�;7G޼)���G��,�Y����{�6[��(S�B��j2��J�vڌ�O`�=8��I�߂f�M`4�ލ�_�� �l�E�G��~��C�W�սw�߇h�]1��GX�Vdñ¹�=ˆ�+��mw�Wg�+���o�U�{.Q��n���x�M�4�/��k�:�J�h4��Ț�׸{�4j�f�F
���N��2�$c���~��)`�C���R�ˢq�K��.�
tA���gI!��f��\f�^�2��9��D�|��܄���-�v~[Q����e�V例ת�fH��K_vrS\���4	9N����Ʌj뷥v��8��E1�3z-�[�#��a�����#q Uq�"t�:�����* ��c �s ��������C�ې��X;�"��C�
�lSNx�͉��vQ�6M�CQB@QdU�
U��5��p�S
4�6K��k�,��4o\jm�����Yr9�K+"����J?��^�Sa���*� i���'��.-�F%]�V��;!���~�;7_�)��/�c I��l_�E�W+��")1������ǘ����k�f������a2�W�H!}V�W����H�[c�&�kuʘ]�hC�e�WO�`ځ���S	�Ǩߣhu�:a�a��.�����Μ��