XlxV64EB    3a22     fe0����XA��_�v<r�;h�y�������2�G�	�qj9��|퉡X�
M�s�����DN:����X��[�u�Ef=Z;�@)]5*i��FS�`ݳpv�ړp��6�����n�ב.���$ѫ�W�1U��j�S�ad�����[N�n��g���N\���[cS�$�(��8A��1�Y�'��Og��,�<�<�"�q���ߵ�JeP���[瓛�$P����袷I��^Oi��~W�n���m�Ѻ���L�8��X2ܬ��Y7�b�Z�pK^��RQ(&�v�IaAkp�M�3�ԢpN�
��c�;'��Cfv�Y��TU�&j�-���諠X���$��z�^��.�B@f��3��lUW��[E���H��6´�wf*��W6�����<c�N��v��L�.����<C�A�J��Ai���[P
��&N�JV�6�N�";;���Y�o�ͺ��N��o$��K�Py�[@~ӝX��"#����R8zۆ��$�v�R�{��%���%���b� ��D�G�P����]��j��F�6�gBq��4�M��,�k �#Q��Ī[�v�k��'�W���3U1C{Y�Z�6{�=���� ���������(��.�6Nt\d88Q�$��Lb���2��G�;���{=bVQ�QJ�������j(P��6w�)���7�@�if�a�ت:�@�o���Wj�J���8������俠j-����jc'��\�
�.�n����e�͢F��\�҂�M����&������_a\9<pA��n7:��t *~�|��"\p-�q�J���G���<eA�!vwK�S3���&���wb&�0,"��X\���A(td�p_�[X_K�'�z<�� 
W��}�'�����Ը~%�SI�a�w�g�9_���0@X
����gB�GSs����e��h�簰$��b�S��H�+!r3gx,�]��lL���L��G7l�F�B���w�&�q�ec@�n"��D�Q�a*;���~x޹�/��*�9N���h�Wd��?����#���6u
Va����.��jf ��=�a렒I�){)drJ�Rz���rS�eM�ʇ�aF�� 2�[���U�]���/��FG����\�����SUM��*a����)��҃����� ����;Y�Li�B��l�*��j7(�W��~zP�qD�Bs���Gџv��|��؂�M�DJ2cs�[������x������?��&j�3�l�u���yݽ�;s=��|�Ou���+S=�p1��'�������|�Z�_�� �s���
e��ہy�dT=�j�aG�H3^>>
 ,x���X����"�]�2�X�)��sC�!,h_Pj=�&��r���)�/�+N�iLɦ@#�硌�}��;�P)ǵ���̤��XV���Z��)#�{����X({߷�H��=��wۡ������� ]�v�Z4�ى��)NF�����!�ig��d6�@B[�i�Y�P��ZkSfQq�3����rg���#�?Z��>��j��-@�a� ��ސ{�\�(�s>�K�����l.Qഴ?���riηD�}��CAV�4+�����u8����2�/m�/�|U�5���ov���T�h߽��B�L+VJ�>�ݿ���e{w�������6Eus��t��9�r��Lme��1�ҙ�< -k������lc�.L$��� ����K�1�XP9�������m�0}����7�F!=|�.�vs�N"��u:4*���=o�>٩֝�wS*-yhb۔�<�&�_�L6��`U\��rq��bS�2܄Z�,��ӳ�	�5���&�x�y���mV�%� ��-9�
���3J�6��!|��5�=�MW���|Ǒܫ�H
yR�޿>���1�r�zPb�� $�����>L�r�H�e8�T�e �MTA���9
��l��UX��T�	�T���&hּ[�y]ɘ�9�ņI�����m�x[`��B���e�X�50(����=�
�	\�/t/!旔�$F���f�v��L�=-�SE֙ ���#}�7Fz1T�G������g�^P�y���D5�����! �$�x�����8'�?�a�cM��H`^nD�a���H8�;����l��K>h8�V��������^$K�G"^�tԪ�
a82���[7�(��x�l����^�6jAAF��5-��PR�/K����������Tq��[d$�0��z<B4?`�B�*�={f/���{�Z/��m��[�ڼ>��=���3���P�ݼ�3*��_D�K�R�e�S���V_�x�����e	$v�}"�ؗF����G��Ƴ+7�@���b��*�͕u=�&��﵏(V�l�Л�=�C�hK�n9�����}9g,�oGwB�b��B��N
_�&�J��N�2��3�B� _�K�9�F�eJ�*��.g�;G��������K-��� k�zl> �j����72��֊�G�h)�`�+���R[{o�Cnj���16����x��E���;��^3�~7 �DA��̻����|�RO շ���`Gt� I�%�\���`&�F!���s�u��K��q��QőG˽�s�]�Ɗ�p2e�mE���^��������t���n�9\��;B�HOD!|�<աXCQX�eT��\Vs����l�w�e�H�L��5��[���P��F������||�T��O�`L��F^���1�:�?/x�G�����n��X�F��> ��IHh���4A�����Α��G����r9��2������RDC��?�$�+��im�H���������9.Q���Y��u�1�<蝭-N���XE���^7���z5y-7���������1n���Y:44��ў�̠,U�}�[q�dې�b4���֦�BL��Q c�^M���hQ�>���
P:�Tb�)�B�9@c����F����O�Lvi�A���Em~���-ث����Ʋ�m��2�ɿ�#i,F�$'�m�p+Q�jGھ{�P|ֱp����#�;L�@�J`��}H���"��]>Ϝ��C�n��(8��ﻌ�=sG��l&���M����1�{@�;�<��3W��8M���w��/.�8��n�J I��b��V���]Of���/GO������8>�MD��ő��pkq�k9'D,��Ϲa�&N*)�9�eUhF'��ɬTG���5��x�Ň�o���8���Q �}w[8%
��1�i�~�~	�<�Lً+��ݦo��E�9|o*���74Y��T+�oEH�V�G{�a-����7v8"kL��	�Wu&��֠Xar�'i�͟yKw��/c�����g	iC�6  ��:��Ä%&fE���Kb���??M��t���[��?�I�6�"@���P%��-���{n��C2��#͕U|u�����œs�.�$�k��H���v.v�H��$����#�*z�4�Y~�C�V���i#�'�7aϟ��=�_�ڳ�\݊:kU��mz�q��r��#PQr��n	V��b:dM:�_��Ԙ�����&ؑ�ҺFт�x���R�� 	BO,L����i����i�dՖw7z���]��
�N��9I���}	Pe]�&�ʞ��g�w��v{����H���jdQt%nSH�#�W`�;
�����S�\�S���8-�(���E0�G�-]�)���� [�S�����+P�]���c�hZ�'���ʇ=
�x��w�
�(q�X��v��I��{�%ގ�W��oM�ڒ�ޭ����l'
�ZK��?�G��
��Y�x��fS���wr����)�Ok<���˗�楙O	���6H���K�D���xQ��}��S%Y�$�Hr�t�jF�L�r0��]x�����=ֳӰ��'_�o]�!���8�RU�����<@��,�����c)M4�cl�M���'7�fTE&y藐