XlxV64EB    5652    1390 �����$w����Uv�����4�{�j��ڬ4JW�z>vd�&Qw1�h�I/�)�P�g����i��5�N�zzN�]C6Q)�Yj�i�!��G@�����,��']�����QMP��N�8���Q����ӂ������u���']@;m6���\�|�~}+��<�6��@�_[�.r�W.� '�I�S��[�u��;��Pׅ3M�pv2A�Xm<��FJ�mEz0	�̷�9*R(�[�+�@p����@��h�{oS��D���E7n�z�� �1�%�P1��2�j����g��λ0�F��%�����ǀ)h���H�Uw��R�t6>���w��m.�0��������⳴q���:3����A��{ISXx<�C�lT��� ^>R����=}%�=C��r�dr�� �_�������� ]�J�T�nQ���q�EO_P�{ 4�k����)UdX:0˽�+`zN�w"�Nan�B�#��
Q���&���e��`\��Qa���fa|�n%/�A����d#˥�Yb����UwZݷʨ��\ N�i03�����;N�����<9^nG�M�1��3 �#=4�tD�S�(/\�顰5��m}Ϧ],Wv��0�ÿ�6�#s9��tɢril�%3���@�H��G�>���ռo��h�]���x�[��l�47<h�@�1���5�d�6��}=-�<8n�aȏPvM2:�R�/���Ec��aဥ�:D:���G+Y�hj��� �8�q̽�&?��e��6��T�-i:N��o?�r�V'�ޅ>b��?EG̈́�U���EQV���g&��C�^Bj����jM����W��������Kb���(�i����W��h�/Y�:ZcG�m��0��;F��?����#��p������G�>�p��\^�mT��y��GݷΜ�	��N	!g~�.}�m:�ڤ�&G����:���9	?`�d8KB5n��-�o4}�5��͕Oqq�2������
&��������.(Sh�8�:k �	��e�ԉ�����ȸ}ۏ��}Yŉ͓�|\��d"��b�ٿ���,@��헇f��Wl�$$��'��2����G�����2(��Ө��,m��{mU�+�3Ǖ��pP��������7g�Jj:`�����j~�:���R##�$�o���}{棞����7���Z(i"�1/�eG�K.�����(��s���t%�{Yճ ��O0��:�RY����:~{z�þ��|�!R�WPm-���s�y¼.�ݚm��H0��_]��an07ɻ����?2:�zn�Y�"���4��O;���F�<L0��~�m����)߇��M�@
оs�,�J '�!Ty��yd�GW��e�]�dՃ���ϫ
䕯�8$BY8Ϥ�%�(o2�Q�j���u:(E:��x���)��F�:g�~:��y@��O�3��Kz,4��S��M��:M�&~_X:��}<E2t�k�*�ڑ5$M� 1}�X䅐�#����S���U��E
Z�����:�o�����&U� |:1�Q0Lw)x��-s(&}�A��1�ah2�A3�^��_N��x_Ss�� �� r(��L�BX��X�2�@�ߢQ���H�V`TO�A��S��Lļ� i����B`<���av�m�ـ�� �@�o�̒x(U�&sh?�|�NUM��Y�T��z��f�ue�z�}�&�Ĵ��hC��`Ɇ�G�cHk�RW�o�l,n�'�����	k���/��e-XJP�3����/��;��U9�a|7&�qf!�Br�����W��Ѿ�ee+�����aC�CzO��YO�DW1{�c�/�>+��1�F�����>��0���N�Zg
SF�g���9g&-�L�� 3�G��zv��?7�s)z�8;˨d3y�d.�N�l}�A
ߚNuV� ��i@^���)ŕOhj$���W���e:_+��o���rIޙ~șSG�ۘ�*?�9�n	p�ǌC���~��8�v�����h��u��ftsOsE��RR�e	��:��5�Ƿ�H���Z��E�y�|�Ɍ>�FT��B�L�+P����eZ}WU� 8Jc��,��[���#����[��ON�#e����c��W�@�I�Ͼ�@+�kN�ߖ�|�	sz:J����jې��.?��T%"���/�&OKG���L\��@�FXXYK�7MrDYF[��X�N��#O��w&�9l��Gطf�T�d��ʹ�K=!���s����<r�hJc�q���z�9[�%Wȃ8H/��u�Jq�.  ]��>2U���4#��J�K5��5�BR�z��v���0]k��7��\Uh'���C	���\Xc�WZV�������"k�?�2�G�c��HC��l�;���b;�"6�r>m�q�*Q�+X��	�V
���=k�4. .�yfң�z���G2JZ/Q�u�]�F�Ȉ�����DP�/=�F��b�#T���Í
_U�E�K���sDth�<�8M�����2o���=G�'<55TG-�Fߵ��z�I���Vn_Ð.b�x��u�f���HC
��I�C^�i9жW��
�;M�.��L�y�%"x�E��+&�>�$��A6�zv2!�v��#��b�������Ap켹cU<	�9�xv�Д��P�ʹ?�n�8�����ޞi	ލa}�d�ǽL����-ZN>��5��/�4�t\�E���Z�$��,��T�-Jv�P�T˱�NS!q���{_:p����,l�K��>Z�KX[[5�8�O1d�U��`ڷ��pi�ue鳕���@�
���-b�nƎ�r�%"�����|ܗ�9p�1R5�bSNi����\��SU��)���3�5^C5I����p�C2з��������sP,�Qc�-���X�z�D�;*�Q3�Aߟ�˻�̈́���3	��=�S���m�Pλ/�8�gPF4����+�1����K-қ�9G'��A�M��{@��i@�K�����n����VM�'��]u]@�NA�ĺ�[�g
�����r�3���}0N���dM��^������qg�[r���_V�@Ԝ�"K��Е=f@kH�����ccM�Ԅ!G3�ޗ�L �NAH|�t�rq���}g��EԢ+Sv��E�
T�����/�i���[�'��Mhc��J
��8.����Q�#�<���oN��|{e��{kK���B���P��o�%6 �}
�&^H�=!�LNۛ_LƝ#'��Y��*�1�X㶱���/w�.}q��]�m]-œ����w�u���O*��$4&V櫞5�X�ժ�mot�Y������XL<�V�b�*(��A�?Zl�Uռu��n��WLj<����?wE/�w_.�(^iŧ7 Z�翧��-�M����t�֟b��� ';CW�
���x�i}F�QH#p^�><B���0��,�g�H'&��*��(C�����K�Ro��_�=�)�l�$�2��VҺ{�z�<�{u�TK�"�z�w�� �c;f��t?�=ю��#�T1^-�ֆ�߹��[I�`��+nX���L�ȅE]&Ң���3��C�n��\U_Hy��S��o5Q;�����s�b���Tb�;ByY�^{uN����\��[�P�y{���i�N��KaG��E�23�*�M�@���"�-ȿ�:�r��a�T�$Xf�k�;o��z�,��x��=��Wx���p�b����$).hOEܤ��9�(��&M��{0)��oKI��x���;R���jV8UFf�Zh�%��W����v����D��7M�nh�ϝ;��b܇
�C@�,��*��<�-�K[5~R3�cC���Pk�޼��n��:���x�1+"��M�9��M:�a�^��NPG8�3޲�Tf� w#\5G��pQdpa�b�>���K�aBsm*���w�GVg��/�sK����h���-k�duS@q�m�u⌢����blP��[UF���f�H/G�ޝ�*���E��>� ɵ`���%��4��u{�*�nzAG�@�`e~fT��r1 �ح�	���Vz����'b�Hi�ؿC�����z��L��U�js�����v�(�k�� ����<���CN(��s�(��蕐0`{������1�*��J�\�Q(���D��O��/��L�����郶w���0$���gѺ Y��� "�<�!m̒��*kA�1�=� �eC&�Ii��ڨ�����>�$�6jOyy
-�?�?��ȣS�R�ex���|���m�<���q�knχ7�I�җ�e�#oi�ؚ��v��4o �M:m��b7]�A��i���sTi�{1o�9�X�z�z�}W��{�4��%jk�ۂK���:b�̽�ʋE�|Į=U��H�mQ)�F�X����	i"s����@���p�W��M��iǙ���A���Y�`�!bP�h��
���]�+�ŋ�~��g襯�5��]:ѕ_zuز��������4�|���B5dg��h2�����ˠ���9ɨ �5��{9��vix6/�C�NU��Ű$��9�yQ���˱8�`�	�1����D!^S��Luj���p!���I9��%��݂w�xԨ���:��u����`*��^���ͭ$QX�}�0܎#�<Y��9X������ >P�E�B�k�>�EnUSp۾Ə~��PQ[�IL�޶�g0vk�w����i�+�b�D�*B�x���^{�i�Qgk�Ԇvp�ĥ��i`r|�����۰T�񷵷�4��8����4w-
+dN��f�.,	B�K:y�m(//�z��y,���׿y/�u���(��+�W<�@���S�«��6���+�0�5w:~�h�:��`ő�<"\����w(����^