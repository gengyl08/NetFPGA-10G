XlxV64EB    fa00    2ef0��p���/�X<�sT����U�x�ˢ����퇣� ��)=X�h�����$��Y0OŻ�6�	G���*HS�r��?�|12��"�}�:��D��=�J�Ed�#�QB�@eϣ�5!{�k�.�ܕ�Nu��}l�q)t��{��r��-�t�I�4G����axJ؂�-�ߠx|V.ӯZ.�v�̖�V;T�r9��	�!&W�I��#}s��O�RC�վ�]\	5��d�`h?���[N�Fl���|5��+y��t&�xS�{��p��
H�R#[!B��-�`�:َ	B�(���K�IFr�8xh`D[�զ�)��]j���X�����+D�m�O�^�/���,)z]�o�'KX��M˒�K�|���m#�������[�+þl@�D����+A1Eޡf���X�K���BΘ��^XJo?H#�_�9�L��ܤ�?($d����bV{�������a��s���C�g*V�M(t�@&I��%h�1O�����M���W�ۋ������4SA�{@�km(Q?�6Ƅݛ�����G�q_f^�������b1�8~�%qF�B/�YZ�H��KK�~L %毱�,�^��Y�Y�#��Or5�����8�8vwl6��}�;U,�a�9۷�	���	־R�,��r	���P�����~���O�������ӠF�dއ��:g��Y�<����`70����ΔYD� O��JBT����բ0J}w(<{7����QZQ
	��g��`�l���V6���b�*�e�϶+����|������&7������D�
qfo�[��zL	.��b�㒫����ٰ�������ax���o���u����t�.�/PU�:��{���ܵ��}�i���\ׁެ��<vf������b �	����O�a���Eү3���k��v�w۠���'cd��p�F9p4�֍�J�i�wv��{;�y���-7�e�t���̛����`�m�&&2	-�?̇��7�[��Ke5�m�<�0]KjY�$�`հc~�q�<�h��]#3�2���}�������2ncok����;Qn6�E.R\�
�����.������N<ڰ�u��J��kq|&����r9qj���t�Uj�P��`pM�B\zkPy5�/����!X%Ƴ�Ǭ�_O��B4U����BYm��z��%L҉c�q�Jp	u�0m��|�Ӿ�W�����t@�f�����s�(�]��8�}u|������!��:���$�����v��"c�
�Z��U���L�����	0P6M
�)�X<G��=L�!���v���j#J��e�{d�w�-�Dq��SwY,��h��]����J�n�F&��md�a�|з3�;�����/T�]d��O�\� �S5��Ȕc����l��l^<:�	�;z�L F��u	&��������"PYKj�ݺ�^��8'/b��-������7�jl^S���:��=�X���-�&�k�%�L"Gp�RʘB�J��-��]���U�i�o��_I�	ES���U�7��8��!#Z�M3V��C8��#�/�%R��cEu�_�e��@��;St�Dw�����S���(�:~~Ӧui�MF���R��C������X�zHF��Zw?�n��p� ����ǏD�@$�]���v�˛Pjq��P�6?�+����m~c�g���;飬��M,�u��ԇH�s�Iru͚�w�!~)7�\��s���Lk��7RpLS��̻���j���{A��z @���{ c�y�e}�Sy���p��$��	3y�v�,c��>K7k�.+�[�xu��W%?/��s�S,���5�㟺�T���aO��t�[��p"X
�
��K��]�������%/aӁ0���`���D���Fs��,��A��K
[�\׍�В�⻁�6���'P�B�E�]h4˭p2�^�,���e����"S�zC7pV+?I����9j�,��"�w�æ� 7���<�]o-�xZ�K{;��q�m�Q�l��>�2���C��P�I����6���\����?]�!�4F�&��vuy�L^Q\��7�s�ˁ�2����l1�U�ap�ke�SEI\�1("�����t!��Tg��Բ]��c��Jw� �w�Ʈ/�h��i@���~"T��o�SE���pNu慉�#f^��a6U������"�w*a=ʶP�a,Vgz�"��H���營"ىV���S.6�>Z.�Tt$�Zp����=�g�I���M!�K��ۥ�;�w�7�ٜ�Zr�呜X�2������ ރ��������
�-��|շe(m9y�+m�Kl�ru:�nk�о�1.�O����z+��ٽp�r����#%
��_j��*z���mh5�����Z�ٸ�Q���,u���_2�cZGi��lV���eKU��w�~��������.Z�� �Mv��'\95�P�_5o#(O�c�����2�ڍ����Hy9��H�L����5:�r��]�s4��޺�L�Ǳl�#�E�ࢲ�l��d��9b� ����qQ�˳�̧���`�3��{��x9iCߑw1��]F���a�7Pbv�H>�2�T[�����5BN�ҜB��P����x'�ܼ�g
��������չ���J� �b���������+[�r���M�-~鰨�s�S=B(�)��{`�c��a��^�'�t;�-�ؒ�O�>/���3?�>��Z.Y�S���o����L$P@W�����aܦ����",�͆�ܐ:#��G��[Hc��?�8l�P/�^���|>�f.��!hdgGp�G3���dS��rI:ɯ�rq�J9��Z���f����%�Q��%3-!�Z��'������c3�J�}�hߨ*9�{~�"~������>�L�W*�"��6w:��-��~�p�'�:������ A�X�����u-�"1���l��.F�	H���B$82�"洬���I��O}s����jK�9�h��|��|�����,�w����M� `��^��b�`<}_��]�`:��\�	��9-�*j;
ٽ;�0���r��>�7f^��j�T��-ʛD��s�ׄ�B�d8Z�
~h�4�M&�-���=��K!@��
�OĢW�q�s$��SK���ͯ���^�v~�]9=��Q��r��˞K����,F���ߙ�Q��VF�I�7{v���zϻP�� �$ �xxn���r�{�������3���4�eg38�s����j�O/\�U�4���fw}�r��QTd�}a����7�#Q@��;'f|f2��V��N!����!��ýF�"������ɇ�?z��M�m>��{ȯ��
��}u�6�T�3i@�2ד���my����	�/# Tf�T*vr&��
�� �UZcw>7Q��IW��i��{J�A�I=n��E׶?S������֩ᙶA_)u�G�.���a)c��ׇv����U�I�t|R��̀���r\�T-{״�����L���4RT婭B�̪A��Y�܉��o
q��z��lv-25��%�Y�P_�ˌ�)~U��z],��)ͭآ6|�w���_y7�NGF�d����f���?�i\�<�NK��_Wk��Rvユ�����{�Y@��h�h8L�fj�vgR�1;L�A�� ��2�<�cqK.�,00Pzs�+˟'�g%����HkrqD���=����˛8���f�;F�;	�Q:T,O�eO5t��)>%�����f��:j'��͉��9V��%��i(U��2q���?���KkCH��������5p��J}	Y)w儖.AQ��l��W�������X�վC��$�
���Z?�R�'F���Ԥq�������n��^�v��\Y ���?�8-st;�m�:V�*=ìa�V� ��B���?��ݏ��A8�c�ȶ�m�Dm���#��o>�;�M/�A.8������m�B|�U�ѹ�D�����SB%Ѷ�zύ��&;m�J�}�5�l�(8h�Uy�|ն��^k8�=�RA�����:U�y��jd��= YL����&DE�`+�L��� �Z}C`�e��U���렃����r_K,fw�W0jWJA�i���<�x#f ��HU�/�ڈg�!���d�!�I=����]��m	�h�8���]���� �v;~�)�QV�8��?J<Ik��H�m}�8$�	C��_�$������l��i��g�[�d�m�C|�?u_�վ*r��$>]�t�e��k��\1���\$t��\��P�򾣜�(/��+�~1�r� �,�[�{����)�,^)ُ/�b�^i��i8�.[E�%�rF�����|���=��N�r��>��!�L4������f��Є��4Ȓ�w��{c��V�b���`ּ.�Q��j�F��Ƽb�*�[k?���1��1������bH�hK���Vó
t�l�k�_��eV�7�ZF%��='j���a�,pw�j:#L��R��2v'g��o~����+$���bj�G�C�1ޙ�w�Q:������CQ��I��U�L�6��x���a#b4�x����E�C��Ӯ�e�o��-{��gUz8���>R&n��Q�S=���9Z�=��>�A-D�ܗ��7��^�7�~�ՋG��{�ͮK�=�nF�<S鏄�R��uQ��˾P�.�:�x}����5Iq��l���9!�㡡�䊴������K柭,���Mm���א�|^�'٫ܗ�TI�p�����q��H��l�1��q?i�ϭ�+�7s�t�F���iMf�E��B�� ��^�}sz'���)u`��^��B�s\˰�.��@}޴��,�]WU�`Q���|��<!��:S�[� �erW:�I���I�d�!B˜��(	����`���
��M����;����?�i~R�u�*�XBQ�Eb�b4HW���{���+|l�*���6[D�8w.ڄ�J�b_(�"��b�G�q?c�zկ&
X0���L�/������V)�r̭'�pw��ǰ�(�@���&YT����S'8�1zKe��eU�+�+VM�.u�u�1|^:�Dg.�< aA�[�Q�1ݞk��!�XƩ�'���m3~��fӟt���w���y��!%q$��~kb��W �[�S��v��z~���V�{{�`�0�b�:Hv�^�$������:����
�3F쮳W�s��Ʌ������ٚ�����c�"uN�*�褉Ҟ=� 
o=��0|N�����ʟ�?���ב� VkP�|���q�`�^�ߦ �TH�7�bl���!�b�N�Mـ^R�<w��p���0#(��<�{��Ɠd�,-�R\�
A9��-��[I�AZ���u�i����)�3�t�m@��*!��AT24ӼB�}L���ӣʪCQ��ȑ� �����2�\u67� �4�m��;�H�PMM׳����8S����6$]�Zܐ��s��h�h]��_ 3�R@�Χk���~\BA����&kR��� C�k���#��AZ��i����e���|��o��/�S��v��[5�[mc������kU%Y{i���\)}�/�ʺ�&��L����)�jW�Q�+4��n(V36@�!Q>�T���O�+�t�"���z�=L+�TQ�V�T��Ԩb*M<��A�텊�/>+��*?��]DY�88���fs&���
��4�����z��X�_V��,G�7�>�u@�+��>T}��/j���BT����Դa�:S�ZQ��N1X��4��F\'J���B���G��I"���/ߑ�h�jGN{�Uw��4�9
��ٽ}�Ԃmd]�Q�"�5�Z#�X�P��8fe�*h�+�|oq3����h��c:n&	ݥ�l��B�Y-�:v�6���\$*��Y���F�C��<.�_3�w�z�Q����.�?n�}�䎇d��c�ħ�6�ޔ�D#B�^ �ƒ�����I_�[%��D%&��x�^:���N6�ј_�O)ˍ�s�ˆ��Dh�Ad�&�"���'�$c�gi�Qo1�1��o�=��bs�uuA�X�*#�u�k�\��OlO_��0;�})(-�*�n�c:ʩy,ĞI�f@5ܺ�SsPAS�� ��Xx*b�y�]��nQ��Bp2��T�&�V�+�a��HSx H���mx�o�G⍩A �t�Jb�V�9
a�W������q-mKo�4����4��X0o~���4�A_�M i��A&�+�􊍅���Qm�������>$F4�v���5v�:�d���43Wl	?Ҳ�2�n�^I��S@�Jf/�d*���l��C�J$2�so��tVC\�a�	���^w��� �E9l��hR�lX�9y!�^Y'���NY�w;&q�\%4�+kB��[�[:����o�%He��{v}l� �G�M*��ŵE������U���:r��F�ӳ���!�BSZT/1�h�%W�pti���:��"]�#���q�(�i=!���l�W���:5�0��[�ꟍ�Q���)A��Mt1��u�#9@$���ڀ�}w����&/�H�V'}w��}<�q������o���fٺ"��k��3��f�h���ԙ6�+����/̲C{?>��g�	,F�Ao)�g�x~��y�K:m/�ѽp墶Td[�r1�!�Q�����@�LEK��i���t�ub1lȊ�mP���Ӥ��b���6x�z�<�v4��1$�G{��δ2W���P}�`f/�O�4�e�vP��� �@�=1?�0[�`�
*�Y[��6�l�� �C(.[��'h�L��w��q_���Aȋ����5)ќ���d��Xv��Q�,#
c��P�w�y��+��]2��o�
5������O|�^ey����T 3���F�Z��,׉��Z�B�>h�����1��
 �`-�r����5��E,�����/�yvP��u��S�@��;�Ԝ�M�V��MM�O�����)����To�mb�E*�l5(ϊ��0&��Jǿ��T�Q7�� �;/չ��"mOz$v"*)�YsE�����yw�HS�X��?��=�+N��)ͩ.���F	J��S�N�������@�>'�y�Žq��qi�~D����,g���(L��l?��ut��zj�wd΍5��Rފ)K��vUXu�v�(}\7�FiS�՘�r�a�5��~���0.3����b�͐DV�xkEr�G�p�<��1�ԂVL��RrP� Ui1IK�Mҹtv�TĎO���rCJоm�Z8�C�����������p܄���f1T
�_�N�,�hq��[�꬇����G?��<�}�%��D^�'\�z�a�m��	'�Yx��BQ3�Why�3�¡����n���}s�E[��9)#J\�N#Ts�g���/�s
�=i
������f;4��K�ؿ`o��jk����l����īyt�(�p�&RP�� ��o6Ŧ�}eHi���6���k��_j��BJoZU���V�*���S P��|�!]l�k����)���d���+��2	��2��ȫO=������7HIB��œ~=��J}݂�|Պ�횜�T���)�6��;P�=��«��\]bI;�e�0TŐ�j�m}�����4��#�˗t��5�>�?}o�!�x�:��Ϟk�J�-׀$c��"�.���$E�Ű��&mP@r��*���iAD5��п����k̦�G{�ƴ�v�x�����҉��y���wN���"�
��4�s)��?"�:p�'���]��*`��b�W�-��	����9k55�W�]]����
�rt�5��[��3ԭa)&KE�L �R��ۯa�	�?��ńؽ�hƣCq�E-L~-�n�6�q��w�/D�cm̡�P����c����Z��u���H�9��T�?��S@�1��ư5�̑$2|�l0)�[Rt����{�	�Im�G����R=~��n�B�T�+l%~J��f�!������Ʉ)6X���7:�j�S#�	���1z�i����oCE�t���f�"�$���?���gd� yuP�wK	1O��ح�����]ũw�\��8G�q��=ԩ�E�Y�I(C\ג"���"kw����G�V�y�r�)�V�G�(>�3UPcS�m�|�����? ,��M7��g�UYW�:�)��[Q�������rԊ+�+D�I��vC0��F1�ў(4o�����u�ǋX|ƿt�)�F���ݞjKbn��]ϰ ���S|�BUxԟ����E���T���"~`�!��O���6:�X��(�%�O�>���T�j^)Ĵ-yMȅۖh�-�@�c��|'�ظ�Vm,������>+�d���U�up��7�!G|i�
���x��hO�D]SZ2�����/��������� �x��~���Ln�V�� J�qI�f��De�m�D�Ĭ�i1��pltIK��)-.~�L�F ��?�/ʹuO�P�x^��t��w�����e�k�R�}V�m]0nf0���;���	wfh��e U�7A�o�p� ���Gn�"K�XtE�����׋����gN֐�F�v�88��v���4Ɇbl��;��~�f��7Y��]���6�
5xR��XC�^��+S:I�-5��LF�s8k���x�t@�v�
5���1��#�,�E��d@���t;(P!�� ��~`��m�eZ��(�
����x�J����6	�3�T�|�s�n� 3�ߧ��]6l{����^�� S����N������T���y@v&T���a�8��h'�յ��iU,1%�rM^���&�"���3���0P���)D���Y�ʗi���"�Wbׄ����Ŏ���F��;䍸�hW���r|`U�S�s�s�ڛ�&�_�w���]�2hu�}ʶ[�u�mM܍X1�5�kHxs�y�SD�6>KK-����b�A��c�	�2�9�K;c�A ��F<J[_����Q�F!�7
H�9L��G���8|�⛍�StZ�8��;_՛�SO@��R��k
��5���`���^�ڠ�ai��'�c�jʄ5�c1?ٌ���b4L��^��k�NVύ^O�N���=\K;��#�}�I�"H�xzZ����F�����ʹ�?R�'�V휩b)���Tջ>�k��3
�	��K����=/0�w�-:�{LD�5�l���A����;%���.Zueyn���p�}��P��89'_�v�ߏ����y%"���rn�K$c�/�55���z����Lv�֡U'	s*�}&��Fj�I��#o�K�V��tl_�X���k�-�/�4�lp1��3�C� ��G7�����X^w��lamC��jE(�@K���{0�h=��������*Io�sڱ�Sh�;����ߐ���G�U�UV���
.ꌿL=���P4~gvɩ�P�� �\\x�e�ތ*ې,ʿ�4T*|�d��1(��kh�ڰ�,�r��?���;�n�,��q�$k!@����i�����mś N}E^��R���bcPƋ���{�[�A�Ǝ�pۥЃD�����C ��,G�l:�1]�~Kn�a�C	5&�!�b0��*��D�N��!p�ѝJ˼��r&�ډ����g��ƴ���_�a�!ڎ�v�U+�~?�mۖS]��.)�׫��N�*Mjl%��p�����н@�c�
�Dr��Q܀`�Hr7�9��y�d�h�|�2.P3�{^��S�
{������&5��$wĦm${3��鞧�(M�_y�jw�C��-��	[w3R�T��{��ְmܿeGJ����p�Vq������r�ӹ�'����Y�q���ea�^A
d�����X�B_�� 8�-"���W2��C�����x���|��*m�y���.���Z1���>�
�@+"'��D�(y07
1F3���< XiS�%<���<������ zH����*C����l�j�ӣG�"�Q����ف��z(?��W���(K�����%f[L�m�W��1B�v���5g6������ӏ��}o���#]���0USz^%ו!�	ٍ������z-�t��_��ѹ��=�,�J�l4�w�Gѱ~��0�_:T��g�(/��! ֱ�l<<,������:�qkn�kiVl嬨�շrC,���nC��?�a��=k{�p�JP(_"8NH�-r�d���1ԕ;��W噢G��9��[����՚c�)y�YQ�W�Z���"N�t��)��֩^B2� ��|ǜ �{a�񻣪S��|��^�yp�Q6�`mC� �c�6і�#l���c(a_�JF��0s�\s`����^���,z*���Ɉ^w%Eev#�@8w�B{f����h����/vGcéi�Hv�l#����\|�d�d��������u�n	Pt�t��R�C��ry�R�;�?���Q�9�s���E"�P��_b�+b���;��_Ūc�e�I�{�����}=ޅņ�2S�l�pE[ǳwY�R�b��Q�������(x�?%`�%�[��%��Qt��T����Q ?�OD#��Zբ 7)�i,��Rm�?@fL�V���d	��d�=�?A�VN�2{���i�� ~��9�p0��,�'A�Kl���mx/Ƕc���r��OIr於88�
͆�<�� ��s��,�O�����V��(���B`��X�2W=�i���l�q.��~��O��}��,����	  �6����p\C-����k��\�+oo0V���:s�����^�	vv)��ȿQơ�;��{��0��~V� aa̎�,��y�E:=
��.���}����⃾��.�u\B\���o6{�m����sp�i[Ql=S=�O\$��^z&�I����*�Ҭ��q��4�����P��8dfh���b��!�f�1��,O�l�/T�Q�
`;����=�!N���~1���2n�"��@I�jl��������>���|�؝C_��r6-FC@-nW,���c����a�!J]E��#�>���Y��e��i/
w�+�'-�~�ƶ-�a�2���B���z�����o$K��*��[o�|5���מ���:��	�7�.���6kf�]�K��悬n8���3 e����À� `�^���L��a8jx���y��j�����T�`/�xY�f����������sg!�w������ۉYb��v��=�ODW�%-u��7qu�η�T�Fl7��H�{=p���8x?��Y3e�v� vNR������Eq�����M�(�4�:��>n��Ku�i�a_<�$}|��m�G�4��Btdc8}j�l���3��%��K����<c�dܗ-�a�o@n�큛��M ���x}�P_�$��Q�"�N���+҇������m0f�ҋ�Y��կ`�Xo,��2����>��8-�"�p+������d<C��w�S((�ӎbЂ���_����d�\��Iվ��Wv���'��Ģ:���`���U���)�[�EJ3�v�Ӏ+�x�<����d#�9ao�+,�ג�s��6iR��{%|)0�O=�h���)�5�iړC���g�/�S���v��WW��'k���y�H���z����P.n$?V�@�������ۏη]w)�C��)>9�`��$PM�|}�f�_�!Z�}|H�<���#���nҧ�:2��I^>�~8�'_�}^�G�rf����q�H+u_�|)��1kKg>y��p���>)�:l�&Ϧ)9clXr��<����ΐ�c�5�c��X�Ík@������M:nQ�y���c94���X,��&�:k�90�z1��_�Fx�lXlxV64EB    fa00    2970#	Ҵ�j�����L9��Tx�#S�8��lѾY�m��7�ߓ�����bi8cØ�?�r��W���l��daP�I3Xy^?{����6�����݅����s��7*��gҎ)���G�C�D�(@ܵ�7g���|J�%��W�x��i�4�q{�`��w�m�C�����@��]�O����@1˒��#S6!��?0�cT(���u&X�a��wϧ���Ѩ�qx����K��2l�=gGN`5�1;H�6@<�?�jw@�������Pt�(�Tn���%h�a�Nkڹ�D|F�Jǅv�a�]���_�o<�����eF��C���_e-��s�7��QU�|�E
Y��E���d�i��m���&��a�g�5�Ŷ����<��yaz�6�m��δZi��K�\Z�
���q�*��{}��)Zu�q��^)��?��K8�y�C�o��^Ɗ�N�~&h�������]sB��}ElZ؃��G��͚�eg̢���ML����`(qw;@-�s�K��R`*;Af&:ԠB�� n�>SJ�X��:�}����.~5�%%�B4G���V �߉ϸO�'���d��o4����x�\�[�s�@�N+��}֥�6�G��$��9޲W�4n�
��`U��� ym9n�w����v ���6 "�T��n��?���:�V�C|�-����jO�Dn���	n����"n���k�R�o��$��Bx-!�8_�Yΐ��ۋh��2� �(��~�|����a�v����	?w
b$�7�`�{��v煘\U�
l�^KM Dh����w��h2�?&��et )+Z�`O%�ymg���Ǟ#��Ċ�U~�����P:{2.���c,�A[E琍T�*�!���rXt`��]�%y�&�i�h�Zx��H?�]t
|�M~�͎�#�*%^��A(W���g�sh	P��}�٪�����8�%I��*�� zOBv��"�Y<|����Uf{��I::���wu���������%D��}9L��q��(�z����������L�`�7��?Z�y��kV0���i-����!�.]�����͔ǡ�5T���'� ��k�G�(,��L'��R��]���s=Bu��@卻���}�'�l��ҝ�|��vƯ��hQ���k���"����7H������ЮEѲ�#E�#�����u��R����\KP�F+F~��:�KA��;��g����@ZОy�� ����)_ˁ��o*�2a�=��2��>��Ѵ[۫�Z�]Xu9�=��<�)���>^� ��L:�.z�4�4�A�r�����U�8W�Es����;XmA�^�Il,�U�T�ߎ��l��L��Ĝ�+#>pPU��D��6n-Ϋ�k!]+��-2��5h�����d7݃B��Q�F����M�1�.D�z�e�.�WR��M�n���'��j�rf3r a_�9��M^'�z��T��Vxm�5����A�a���Ʈ��8�w"�������*�^Ѻ�S$�n���@h��B����m���5��̐�gy���3�x������8d�񛩐�v��-��%e���+|"����(��X���/!QkҎ��P'?�n7�BW�	�;�mg<�V�C�Dy���WaK�[�n����{k	���m"i>�����O�,���$@v���Ou� �S^ŸxA��aS���LLX���w��Lf�����U��h� �|�LS3$Z!�]I[�i*~�j�1+��z���,Zˏ^����mL�����,f`�*̊��ȧC�d���;�W��z�^^��U��������^��<������Q%{�6�����#3���2�����Ȟ��;#��l���C�Q$��Q��n��Cך

��W�ߓEfK�C瀖��
$�υ�:}_.��1��f�X��{�<A�p6� ����m�"�"��ER��'Y'/xM�Y�ɪ�Q]������SR�)��H�� e�s)�i�H�S�Ȩ��ը�S��c�`t����:��\0����V޺�k�U���-�6�bB��eG�9�ҋ�(�x0S洄��8'?�L��n?2}i�
H��r�d����h�Pxg�~e��J76�i-��& tN�OFv��[��?f�_�@|���O�Z�K���X�ME�ES�B�W\��ڇ���������4@?���%��|b��i��B�o�JO����zkW�d��֮�kZYF'�]3״�ͷ��A�Ѽ=e;Ҹ��3b�}��r���R�s��L�A�._��괧�o�n�%h���:P9��M IW�3�N�]�u�V(g��!�!D��������0�Ĕ�ǥ=.3K�~f7Ѳh��D�S�%_���2g*!�������~H��:�i�B�-u�/a��1���h#iI #�9�fX&�y��f�_�]n{H�]�5��hp~+���s#��[-x����j�\�>����`�#�tlu�xE��PׯDƑ����D1	U���;�h���:c�_���=Y�q��&}S*���!�#BQJ7�S#�k8�Sy��$~Q�۶YF�ܩ�<=�>Ӕ�|<�<As�`N��1w"8G?�_�M+�}�6|#_H��7�,��Og�$��
_?��v�D;_�t���HMBF��&y�_|`R7��@��J��+�	��]J�/53�-ws�י�h>������� {z���Ls���nw Y�؃2x�� <��%8��b��/���貜�׷�����<���ÃW~��v��j��u�����mJ!q����Q��<K�n��)��l�C�������0o�r��cѺ�N4I�!��V�o��=ӈB;k�%��޲z*;��!���ypl޻��zўr*O՘�\v�5XT!��W7�vzD6L����P�a�Z\��rp��=����M^������t�U�ˏ��4t�~(8B0�������zG�z��l��]R���{����t��KPd�p��@�'�I�%WJ���,-�|��
�=n0��Y���������|l�L�#���% r�	��Y��I�a�8�H���372�|��z�M*o�'׹=�43���"ԯ�[�Ż���摏��ྼBzX[ u5�%���C��<����aj��[�
ݫU�N	[����+����?=QJĿ۵�U��Y�Ͳ��R����G[$<��7K�(��݅$�T��y���� ��݃����fg�O���JL&���P&��9u-I|�ug��0Q�G`�������n�+^���k��{kԵC��N����)]�xTv!/a99�6H{؎\o�~��_q�تX,���{n��~�~^�:Q|�Q��6��F?˶�4�<.����>o|��N���O�bj�Y|����T-��J��Oh�P#Ӿ�k �AX�߲�:�hP��N����iL�/��<UV*���+?�0�a�����g�,�x���Ϻ��0��ۓ��H��"�l*`�����œ �$�2<�Q�,Fc	)�`BYD=���iˤ/��4.�8�K29�+Ř���d�h����Ћ�QǌG���qK��>V�{��I<_�#���d�B�v�(�6�iEDs��s��~U:W�����w-S�P���8���X��V��d�#�f�O��<}�_��	\;�ɤ�����r��9[W��K���j{�b�)�JBO���/�dAfj*~��M<0).���uq�����V�^]�7�3Mtr� G,���qCM�9ݙ7+cn�8ˆ����gIkM���j#[���r8�J���	*��M��������^���":��{-L2�&f���v�7L��N�E���txq�~ht<�r��W@t�t^=}��K��0�$�͜�#ۀ6!�8_�' �c��esB�@;6�=h�l|[R�(T�/�w(1j!d�N�P�0*;������ܤϷΑ#����{m�����w�\W��Z��u�s��"4h��'��m�^00v�K���s�V�	���kʃ�[d�h��_M���4o�d~��.�	n��&|�;���c�K� ae�^zl�D���Qˏ��!�g�9�}�@�,v��&{	�a�̳�
(�^K˷P�f�TS]�,���9���Ԋ �8��2���rߥ���͑�;�(S�Vo���G���N��9[QÓ1mٜ��y�MdO�)w+��1&m��??Y(�Iy�����]�]����m��o&]4Ki�[i�v���'����ǏE�j�w������.�߼[Z1�H�z@
�})�ۘ/Tt뙮۩/ϧ� �,i1ѣ���K3�o�Ůw2���(~~|X��Wv��~C'�X-˙
q�"㳖E�@�$�6
Q7�9�Ȓ��~Ԟ�<��BK����bw�ǌV��]Tjq�J�1�Ot�344BwQ�|9�Ғ5�Qk&ɾ��1a�
���\�)ׅc��@�{3"5.&�$�����p^S*��Ҳ��9[9��iK
Y�,��7�l�Mze꯽��V�!T ]& 2C�J`��E�K����'�l�w�:o�j�A����F��;�L���G�aݏN���A_�w��r�B�V]D�Qd��/ \�jNd\<�	��r�V���xp��-�(�X?ev7q��W��b�ڲ��w��1��Q
P������L�^�$*�0���r</T$���g��T}qx��g�?rIC�'�7avG�2��YNh<���)7�7�Xy� ��W���WU�� B�Q��>�b"Vj˵���PM��w1D��V�^�4�2�ǭiD!�S�fo4��,,�:*�iT�%X��^��,�ҋt^�H���̻�q_7Oq����>�^M9�c3+�\C���8N1����I���'|�ư�9����y3���nU�U����F�ʕ;��(�3����E�4&�_DH��s;�����.�L�IC�+g�!C����(K�4�VT����~0w�-p�f����Y�6 ���q�>��AW(9e
b��+��G�͇ Q��`|j�
�tJ�6���!`w5���,9�X��ńB~��8i& GR7`��s%�:�~/�H �T��9�6����\�d,ŏl�h /�um�)ֺL��o�ֻ�����>�6��i���ve��������@����Ӄ�܅�w2�������ҽNb����Fe��~�$t|��m�Z�a&O0?��Q8�����9��������XG�?�U��҄�����G�i�k�.�P��=I�/�с�{�T�ŷ\�l"�.�uH���u��WY��/)Cv �&@k�8�Xk�>�a\�T��n�Q�D�LE(E��CsxF
.�aF�HW{(l��Y��(�P�Q��t�s�aU�tL�cUn�]�9a�d��v�Ԣ]@$�n�BL�I6,��Є�I������!	���lR-o�R�7D	ш��DPTv8�l�D2��0t�)��]ߪ�ևGn�qlu���L�?�Q��č�ޞc>_)�m��w�]C0��+��P����T������ K�[�\�-��e�N����M/E��wQ*�4����H�>�Č��B��Ae����K>�ɞ����௖q�CQ��L9�k�ƒj��tW���+isq��)E�:m��a##����9gJ�����r����[(���c�
Ͽ�5-�#��N�.�7�vH��Y,�ޜœQ)u�&�I�������*QX����%E�����K=7�v0�������pO��<����	�_�����N�-us)^���]�಍���6���]� �~��8��ҕP㌠,�_O�9s:(|yf��V'>�!v;%�%v��V��"gx#o���F-/Gx�LH& L����٭E坃$�P��DEZ�������h��\��I8��eh"V��>�ӡ<_�*Z� �]�<M�f��{�d�3������P��8����8��9t�ƶ5_�as���dQ��,n�)yp��D����a�*�7.�3˽���'t�5��I'?ʎ7֢��_�ă��D�T�.X$�1��BZ�����a�j��Q�����u*����\D�=J��^[3'!�3���ƙ���<N���]:WH�u]7pw0�6��A� �����[0�:IuɦI9f��gr��G\9�	Zc]��	H�z~�������0H�����	.���^�گ��+��N�oZ���l���E�y�ĭ��L�^V��i��]�G�8�E�Փ����49 7�=��t*z=�7�������"�,`�˾��b{�6��)��4����D�S�7����U5� d��] U ��y��h4��Y���N��䬑����H�e�@��u���	�:�¯�F4�L�,;��Ӣ��q#I+�V�ߖ鉜,i�S.��>���)�Pmkk����~��q$��3To�k.(��c�r�xlJ�|��b�0�'�tۺ��+ֺ��jP䀞���|�H���p�n�"�)��1ɟC[z�U�y�b�&�[$X4���$p�;SznmD���AG<�dx�]�,��m�A�ٗ,:��^�؁��˷�?�Z+�c�Ԙ�4��2���Z.��Ib��?�0=��L�Fc�%���CS+驉�I�i��X�3�4sT,�pl"��2��eآ��\%���`�����M��GG`�\'���8|�k-�_:����0�z��%!�����$\�q��_(�x?�sC����*@��sWٷ^�Ai5pS��-^p�'*+a�M������K`��;�}�J���[��7ѹo����q��˹$���/ g��^���
3�?|��g��vw5oq��A^1�2��iø�ďp�W�q.f�M^��a[1��{5VX��q���,�?�/��L�m�"T�W�V-I�;wY����*(����z��&H�LJ�F*[c�t�3Q�p݀���9�����7���B�e�!,�"����ݶ�� +ua{�P@_�����R���¦<���r���x��j��|rlz�9��x,Y1�˼��𧴳��~���'� $���4�������x�e��s=/�N��7�,a�׮NB��5��\5��%C�����Ҫ���L��p�vn3�k����'/���a���T���VV.!�t����镡�Җ�/�;
"��e,e&4FoI%FG�^�OD0�B9?{�:��x���_�j��בz���!M#�cA�4�x�2�KU�$�u�����b{��:(e�@O�o��7���(���b���L�'�=�=3v�޵�jE9�he!�wD��~:{Π����6x�g�5÷��W���\�;�l�f�SS�� $��q���?	�[e�`���A��{f9��U�o]���d#��u�*���zF�~������������X�~��Ӂ���ql�؜ ��t"�zG�z��u\+�C^����\���P4K+����E� ��5�e3������ v���soS�������)�	36^<\-}:�M�nQ+Sx�0��ܐ��M��۷5Y�!�sV�_�}�Lw� =E�ͻ�a�
_- {v�`���Ŵ��?Gw7���D���֗�������~�p�YI��
*��P@�5n�C���I8�d�۴^��2������]R�3�g����ܖ���qZak(�i�ۓ�_�%�_���Yr�ox��kLDEO��̿^-I�7_�<"�ik<�]J���:�յ�&��[S�$uk�bdAG/�4ìu�s�_c��5���Tf�/�x@T��!���Q��ȰH�i
�
�ɰ9s���' ���3JP��e�w�A�d��C5"E��)������N
��̡ʀXޏ/|���/�xrr38fq;�Qd84����A5��i_*1�ԓ�]`Q�bY�V��9��ƽ_��(i{pF��аw�d*D�Tqմx'MYc	��Ԏ�d�%J���$g|�#�qWC;�� ��Mם;�٬#q>��� ՛�Y��"��� ��^��n�A��M��}���w爈 ����*O�ҿ8;G^��[�Q��%�7k���~Jy���n�ڀ��}'+� ���1I2y6 �)�h*	W��	����\��R��f�V�#��jgg��V���e��h=�i(���E�[η���NgE5�*�Z>I�`U/���7a���9$:�Omc���%t�$[���#䰛C�E�Y,�=:=e�3�Qs��ιl��P���u��F�*�«���D�_x��jĒ��� �S�\�4ZEW�
���#�
vG��l (���2<;���hg����#
�C��O��S�o,	�Y6�V&�R5
]d���U}�Z�Ǎ��cي��SEb�[��j�b���_���%�c-���k�"����ƍ�� ��C��X��`<t�"YD@~m����L���}@��� ��X8��Wh���j�����80 |T���k���������������V3�WV��zyPw2��RΈ�D�1ԘV*
P���Bu�S�� $G����Ăj����ze9`��>��9�E��!��O-��U��8���a�}!��= y=�b�#N�#�W��'��8W��+�=W����)6�`6gt/E����vĘ����E��|�=�����Kü�Ȑ䞛7�]�v�eV2B��]�z`#!�m��:-�n�υ��C�M�\}r�Y���2�*���.�{"��~�D��%����Mw8�)"]�	�8��;��
~���͏�(���;�7gCb�&���2�N�O�\��|~V8��z`9�A����l���d'���?-�(��ݢz�E�D��5V���C�fc6`4݁�vPT�����m�?��n7}��q���ҧ��MD3�9��U��Bb�^�Leˮ�PFU��nډ86L�FYV��| 5Uκ���h�� T`�	%�%}����f5�^=t(���{�T<?Jb���|���8�&����4C�?zml�l=UJQ1Xg�
�h���%þ Թ9: ������nh1�[j<�}�����Zݻ��ĞF'ɤ�]���3�O_�St�cG�N���߷�'6oj@(UE�'���6�?�s0�y���yu2E�-6��wRhփ~�'�~�w�q�M�$K�rD�ؾY��a�R-_>EDi��T�&qo�'$�%x{�x(��8#���_f��v��Fh���	)�\�R��[� r��ߒ���`Ze
s �q�G�z���N��}�� ���g�� ��V��[��i��� č;-�[��,}f0S%rDMߣUFgB��w1Gu݀���.�V�A3��W��tZ�i�>T%w�g�������4ŉ�H��	QD��i�;��P8�<�!�W.�:�����J��k�1���*����k��� ��*	s�g��.w�d���M~y��=����=z/fS
c���D*"�yH>�b�t���"�͝�ʖ>?X-�]p U���!�1�rcB荐����Jp��N/H#��h~.&\6�?����eR���:_d�b�6b��nFTyCJ�~m�H�[H\�.A��%����9�K_�
� ���$���������#T�J�v�7VU	�6
�e���M�m��K1D^��GtJ�C��&KU>�u�Y�H4�Œ\����g� �|ˉ��W(e�;�؁M��:��*�Θ�3)>>�d)#<�b��-J�n�l�5� ��c�$����n�Ü�J�D0g�e�TN�f��s9Kb@#Z�r[�^����������Tw��-��
�+�S�B�vN�I��x6t��G�~���j����7�$��zs.���9�O�	%5���"�p4� F�x����1M��# bΰ�h���z�-��}��۴_��BH��`m�����:[K�{�7�E�)��~Y�o�W����ri������cW��p�Y)�lp���Z8��)��#�x��6��l��{���@l��H�o�kS�\���B��5���2��1Aӌ���Z�wк'&-A�YF���}�c^PU,��&n�b?je8!��w���U#h_�p&%�y�9�u`(�v��2P8����%��v=avIqy�Q�����4v�6���l^����^{��Ɲz)��UP�K<N���^��
#��/��)��<�h�������{L��ؘ����{�`.z�f��P������~ZϜ���+	�#����#G�av�1ʄ��re/����|0��R�  ���<E�A���-��M�)��*���Y$��D���z8+�iܺ�,�[l]�QX�xJ�Q#޼kn��$�����XYr���SO��걑6�aF�ɗ����4�_��v%����+�P$KNu�Ҍ�=� �Z_���h��DY4VI�|T)n�v�KiI�B$�!=ҽ@6h�ؖ҄���/�|>9�iz��XlxV64EB    fa00    2a80	p��İx�`��T݂��P�C�#Q���J�/ykA�G��R��-v��Ԝ���2�kf�Kz����׼�q!cT9��d�ǜid`��<E�3��Y����v��G�#��=h��~������t/{p�oh����%�{�O�9� ?
v������R��f�,K�W�'��Ԝ��+�2i���$M;��"2���6��S/dn �/Jӝ���	�D�ÊP��Q�V�I�J����M��Q��4��Gg�B�Cs������x^�okg="��h����4�ᘌ�	�Y$u>ʏ�e��Ѓ`��=p%��T�||]�������ZCl�s�����<ss�Rmh��+e[�h�CG�{� �)@D��^���ꠅl�/����s�LK�ǗQ��A�����`��D[Ω}���GZ�ϭ'����&��E�z���u�q�Y���sz�Yl�Sp��M}m�[%`�0�79�z�hR��G�3ݏ��G".d�r�w���1�l��VHe�rE���?[��|"䜚��k����/<I@�X��x�g�H�E�L�|��ںєs9�C����_C�e�ۥD�ہGPY q���'���._t{wF����Fr.6A�&=�L.?��vyq�\�*x֭�������6��-�����){dO;�RFf[�_�N1�òM��:�҆,��)�V�����X�d�o�����.h��l�Qq�ӫr�avS[�`�C燜[Ge�
`�	��jH-,oH��$������Q�0�t��U��p䦧��:�l�q(��M� ��Vr�� ����h��2^�h2LS&ꛚI���J�"
���������0�?��ڭ�?r�C/]9��H���D�
b��ek�+*��m�YZ@Tx^�X���%�����Ȟ����*;��%������Q��6�������k�%7R�3O�W�9�V�ޫY0�(����� ��P��4a��8�>vt�tz��~oD�J�e�Nj��WA	�f�Ӫ��#S�m�~eH}��]��?i"�I�36�A۬���p|��)d13y1Ҽ͜6�O���A��*+���G4x8>��{f�nD��ň��L�.���Q�@l�C��l���$OlL�RY�2�ȴð�z��-�F�WF���$6�|Gz�gtR�M��i-��`���i��
��Dl0Yy�GXj�C�c�+F@�w꠬C�?��R_���~��^�z�Jp/�%��V��#���=Į���y���;�^9��<�F�t4{����X=au]��c��R��t�ٚ	(��R�<��t�0PM�-��ii��3�fso�4�{N[�BE�𩤆!\,D��_��,�n�:x�Y���8m�cr�̕�P��Y�JQ�TքO��ǋJ�`Wݬ¼�!�@+����K���-|�����@� ���#�9�Xc�m�>̋UNUhBU��p����7�6Vɉ���J ������ r�r^t�F�AC��V,BOC���Z�S��[f_Ո��[�_p��B0F��۳�6����'�S��$qUda�l�M_�q�vm�R&?�qn���J���7n#A]���|#4��/����T��r^���6��w>��G��X�y�Q�]9b�LFPxc��4Ꮌ����z��YqnOt�S�nB���k�`+�Ŏ�:��7�"d�I����UDk�6�R�[gFZ+��]�&ȓF$����
��2�F,�ԚDkh�B�� ������Y4C\�ư\�5���2��d���
�]���E7'�٣ ��a�2p5�Q:����\�Y?	��dG<�y|H����9/�ipݾo��h�d��^���㰛H����Yt0D���� aH��$&�^5���K�*��ӌ�iH|�ݧ}:s̓�*k	,�̆!���!p���D,[$�
0ۧ%�&����s[�ڊ�Bk�i�[�#�GƸe ��z$��y�(��lD�=��\%��W��(le���"w;�!:(+z~����(I�m:E�/h��Ӥ�tDz�`���W�դ����f�4�Nybu�7�{�Ʀ�����b��������-ni�I��7�v�o(�v�����{~�9]Y��ag@�F������_p�:�,	�ԛ�d�m-o�w/R	'd�D�_��FPܲ�b~����� �qL*u:i��'@	F���;�_���Ll|S���&���u�K�:BϤ�^���nё,(�I�><����_uK�4�;��ST�w�b��6�&T D���b�dq��[���S���Z���b�<Hm�pK-} f�e���_hCS͝�cVv��i�L���WܩT��F���$�Hg�P��m���o�Qx/E�e�@�!rY�����"�UA�%���,$�c�@JX�iNUZ���&1P��j�Xxkٯ\�G���vB��Ѐց��0-�$���nr�$*��B;�`�P�����H�J���/ȉ��&Źt�}�q#���%����wu�b(�����Q�|piT�V":`���!�㰂"�5�"շ�!	���tD�I���Y�K-�!��A��cT���O``��P ���F���h�S��/x��bN��+<��gG�y�e�b%������0����_�v���܉�K�z�GY�v1�l0�,�E���uBݳ�_�҅g
NW(��7L�#V*HM\�"_u�N��R|�)�1a��֤ ��1 ����D�
�MO��� ��g�B/��~eJ+�U[�.p�Υ8��$����	�|�����N�v_"���������e�)8��2��n��g<86�_(���j
��L�jc4��?{�܀�����;�Ӫ`�/Zއ�S*�屖j<��{m�C�qЉ>	���ka&�gŷ���J�9�R����l��a?Y-�;�{f�ڤ|��:�8��oOk�o벺����+��9#��{�d��WJ傕���Q��۷Y��������iw�ӸK��G����T��1ƹ��j��#l$�N��k��'KŲe�:�k��-�yK�t45�	]�A<sCd�/
�4P��V<g~�̇H	�j���$�����^󂾐�|�ѕ�Hq����^��٩{E�`��*���h���و����$Qt����	{�����Y���_D��?��aB��7'�a�6����Э��h
m��o��X�t�-���i�u��k����Y��g��"�
IB�b�{����C*����m���ς���ǋ�xy011Rg��R��-��I�[9̸u� "�Y�f�q�(z�U��@��`������+���F%k�Ƶm�a�}�Zv����(gI��3Ј8Vz7��l�t]U�t(V�7�Փ}�^1�w�*�������t
w��[_���I%ҀMb��!���i>'�ͪ�~1�(��n4hn�5Z��E0���)�*�񅹼�Rne��u����
������2h7מ��K���!}�:*2���Jz�]�Dv�<a�\�ϧD���{�N�<e�1�Z�	�t�D��.%����?�_�ι�7dV�L�L%��|Y���WQ�\G�҇�.\o��$�m,��S�UՀٍ]���c�-/wXO � �|�R$ z�T��z���8�����Ҹ�)����8Y�Ǎ��S͑m߯7Mmt��ǜ> �.���N(>�-?,m:�\1��N��"o%�>_)3k��Ni��șMP�GF�]���\w�K��$�W�!4����/�&�i�T���45T���������r_�����SQ|�)4�2>z���!��pX����ND)�>J�(�Ɵ^��IZ���X(2��M��)��W�s��ͥueO�״���x5�N�q����61�zf*��O��,�
�At�q��V�9Z;J�У�Py��\ Gv�|���%���_qgJ,&+�$ґ�-͠��D�Z��"�3'Ys�������q	>
���"q��(�i�괿�����]��ZJ��mQ=W�ET��Ա�τ�E�/����S�NB�_�Z�e�`�j�Š�	��)g�KpD�,_�'�}Þ���c��<�"�'��:VB�sA���5�JA���L>[*3P��=)�Yx��5��~���]�(є���zb���2�oTB�u`͚Wv _I+Se���|�]Iǫ'�3���O�/��k��2�آ�xB��H�wN4��/���s�߅��7s8�p��l���i���C���|+�^�n��qEQ�V�J����-����$-0�V�n��s���gU���d���m:B46�����4}����\�#��#���8��V�����=y�f��G�Xw�����\srbZ%m�U�eF¢_n���blŉύ������dh�'����òj"�4l���I=Bc��N?�d��wY�e�ӖѺvFi��)D'zi���?��}^æ[����{���a[�~
��4��V�-��M
odSŜ�TV�_x�P�C�܏_�ufE�f�n�|�tv>�Arcm�ﷴ]�6ͬ��x�כ����|1�WQ1�qӓޑ ��!�"�uvێy����[�&�Ә�B�S�eJye�/�Vt���Sm���<g����tR�c�iB���{�Rn��@�g	���V�z����p��S�.���+k��kU[+-{�<C����U^�x¹�ɵĲWL��SYj-�8�����>K�hYU�we���<A}F��/�������ƍ!�f%
�b�����+l�2`gw��y�e�9���;�q.�џ�J�E  ŌS&~��=�2�I���r/B�\�[B�|9��C�!�Bx7��<Q%Q\Z��	�ś!*�ߋ���L#�k�h�F��2T-;�
��n�zuB����	q4Q��|Hh�-�פ���6x����b5(�b1-�G���X�ie�Y��(M*I2�9Z����rB[�(�囕�y(�¦	ZM��`#�F���Upg���:�
py1�s�bI�^�V�U�?�rN%�,���o���u;���1:$�#ץ`�
`�,(�\�L�&f�b�x&��a�[-A��1ڪo ���cS���V���KwU�Tc�P�_C/Ú<��ax,��u0�hqC�6(@D8N��c��N���TrO��:���D��+I���E��2�HuR�2�؂bζTJ.z�b����E�veT�1����l"�c�D�k�[#��%���������=)l��u�&.>@��6����YBv�R��6I�e���x/$�,��H�Z���?�Ǯ~�/
���8���'Ԯ���2�I:�����|�l����F��ÜS�su��I)�[N�q����+�MK�d���[�\C�Հp���3�>�z����l��о�2(�?��|�)�|�u�%�����玾T�Aji-�!Lߗ+!1���,D�hp$�c٢�3I�r'q�vٗ�wS��M}���}�f��K퇋V�r~��,��ng�I�c�Ʌ {2�+O�Ag���]�\L� 	�m����~\˜�;
��sm8��k�:;��ל�)5�px�Ӡ�K���K3xP_-F"�Y��v�u1(r2����� ���QK�h��t�ۄ�v��Ɂ���+J&��d��W�аQ��
l^�)��L�.5�M�S�<(��Ը�$شO��m*��^���&�g�m:<�N��y�8�Mi(��9��� a�1+ڠ�3����G/���ѱ�k,����䳁;���wg��&�[�����h�9��	c6�6^j��^�����^�Q�X�N%�z�Q8�C�O�Q��,�hm�K�W���CNf�P�� bx
]�[�_D]`S���O%�Hɟ�F��?xP��gZ>���=#az;��$����3YB %g9~�q/����gus9�}���S�h��3�W{�1�{�p�*?���l:F������eb`�L��=��pzA�'�:6W���r��,ˍ��*��@tURS_�<���c��m����}���8���|#�R]�2����*鵄�=𤋮��·F�J7���O�()>�x��V�Q[Z퇽=�_�� ��<�T��M��p�|�r3>8y(RlG5+] �4wn`K
ͦy/m}������a����~X�l��-wH��2������k�E��aҕ;t�+�Y��`��&�PM	��F;i�P)��.1˒��a	ZBh��Bwj�LUIO�ʶ
�Z�ȍ���Y�|���}�X`�BU��A @�Σ1aை��6i�*���Bi�{$+;�^��.�g�沆��q������WR��_�Z� !��-�D��mD��p�oŬc�8s��g���y�5�5��3 ؤ"T҅ �h��W��z��0�U>4{��S��ޢ׭�kS0
��>=�������Q^yꯖ�L)D4���(�̽�+��-zr8o�h�;E(���d��b��p��ў������,��"�c�����_&���9��i3LQ�fɻ�Y�eL|�$wkhn��Ƙw�9nx�D��м��%��f��%Ϻ���un@IO�HC������W���sRp`,����Y�����j�����p3BWv|�������qȤp"?P����VC0���׽�U��];l�`-������p�C�7 -ɻ��у��G��P�jpb�NQ�k]ଅ{��e�,�~�BA��H�Y�n�R���i(4$��]o����<��v��X��0�/�9�)�Z#�5�T�1�/q��*��>��'x24$nZ�H���t1�>�?�A]n����J�{�o�K+"�����������i�gT�b��u�ѕ\���u+T�d	遻N�&b����~\�x�e��ר�o�~P����N EiW�Rx��ۣ-�h���z�8'�Sԓ� ��#�Uy"
;R��^��a�G�9��
��7�`<;�p�u����l�/oɞr=)�zg�������ܘ`���9�����^�S鱾������WV�D��iJ��s��o�0��'P8� $�$g.R0�Ѡ���������p�9�y��nф�}��b+G��,���w/��ZPp�Q֯+v:�*��ɕ�p���ǲ�[���S~KP���q�w���sf�yp��`p"��f�(���^◻�����y�0i	�o��Z-2DԄ��,��u(�Pv�h$�7o���
�0���6��p�����I Зv�\���ʫ����K��F�
�����!v� O�Oէ3D������*J��;p/� *_�)�ԇ<9��Р�8i1J��%}����o�/ӄ̶���{\�3���rA������S+�2��wu���:�Ae���J-y�|�+{�[A�	�~�P���"�:F�����R��p�.U�sJ�Ќ�X���]�D��M��6��0Y������e)��ܡts�u������@���"5`�m�'�ڲ��u��3��F-�͑�}��E7��^Y}q	f�yJժ&����>��!�c��_CA�#yD�˙�r��|���
{tAtM�Ԝ�Kr+h7+97Ń�rCzw� p�~ny�������X���\���c��y�q��.N{i�ca̉��؞����1���>��(7t�'�f��=���p�3����jVS�^7�'k�'���W1�$�?ē��3����$��x�?�2�O�=�b2���a5�@�Xw�˾(��Ə��`p��J�}��#>��av@�t3�~"��V���粉CK	d��A��y3�"B�e�`��wv	t��eQ�0<v��������8���y['X=��.���.�D:��;�ACS��k=b�u:����bÌTǸߖ$b;�N��A ؒP�2p��F������K�'�da����F�9��n��r�:��e���z�.�X\��"�U��r����<��f��e�K�Ak`K�7�}��t�`j�'>�>Y#�Q|]��knIz���72�J�����s�76�܇���.���v�x��v<���OP����F�ˢ�'z(��u����o��t��e*����󢦪�ڊ^��~W!�$�?|���V���,�'= �������r��+�C_=�:��s��3.Δ�I^o6��^�9�ޜ������raQ����� H��p��\��њ���|&/A0��7$�H��Nz��y�_�g�������ty.17�D��W�i��N؟Z��\,���CcY3���V���k2��1���C����H�9Lk�a�׊\,��zkY��7�o�]
uK?`T�����kw���3y	Kh�߮ʏy�S�mϭ�lb�HޑR/�G�q��]��~�	�°0)��uM";��DCy]XSH�L�:8�����.�5�#-��$��]����U�0��X�+wi���.��4Ik�rl��M�Sj!:��W���g�%�Ƿ	Dv�A���n�(���M�65��1��n�CO���YF�ӣ<���r�+�����fDjQ��qs����n�����ㅍ�s[i;F��aE��x���kdDzEb/א'�j4	{�R��c��CWH6�2fj`��>���b��Q��X�
��sv�b�o:$���x��Jg���|7Z�ISZ��@-W6G�(3\'B��q�"\A�a����1��-S����a+u�B[�/��%����,/Z�1'�y[��wOg2,Ī�6�|H�fu����V�c�i}�&z���s��a��+*�W<��a�=,	��CVb�S���7��(p�����8��y�N��J��o�k�]Xuj}Э�����5���Lỽ�a��s0Ŷ3_�u��-Gs${0Z�V�o45NvH�޼Y���_��y5Z?�杈1|�3���@��>a�������N��LR���v���yZ��� �M��קY�z�ç��f��40�:PU�Κ����P�&�
���l��/w<)� ��Q�t��Ng��锌�����Em>�QB�I�����U6�Q�qiSn�ơ�T�j8�|o�)�֨�����mWƙ�L��q0�i���8c!L_N�R*������6_��^i�'GF`\8��܋O=�2g�z�e=z�,�M��TsWYYC���xw�ds����U��N��_�
�S;=�9%�]1k�E,M�&�����^yh�%C"���B�����^��+���tp�^_z����Y��d���R�R7	��rٻ���%0 ���
G��R쯊��m��'�"�+*�9�kW8=|v���h�s��Dy�T�!C>�?5(���yѐ#�Wj�����,��Ð���׾�+��!�������;�Ҫ��fhP��vf�,�R��ղ|���~���8�ud������Ƽ<����"#n���� ��h���vh��X<�Gpq�2YWr΁��Vi�G!���J�K6B��]�^�^ֹ:hM�R��6��L�{����bÄ�����Q۩�z�z<{���3�LR�С �?�
����T�M�?�o��%Z�#�C���&��: �\����ݾ h�o>����ۦds �K�˔s���x)�d��{�9\2��dv����R�W��'�!�ں���R����T��[��ٟ�I��*Z��/7C�E�E?��y�E��~`�\�< �d�;��1�����L�)>�zk��
�UjA�5�8�<�%p�JXÃg���~��យ�˵��oe�W6�z0D��]̫��{_錮�hv�5͆앾�u���7|Α;��SS��g��6�Z�l��QQ�]��y7
'�Kx`��٨4�w{q�7����-��\�*��J�c�`M���д���w�#��;��Ol�C�=oˮ���&q_E'u+?S�RGt�)9)��f�h-{�(g-�HqW�ck7U�5��o�`eL�8=�B�ᦧ#Tf"�����$G.�xW+j��8u��f���.3�����33���Oa����}f��>�m�k�G�W�g: ��o�KXc��yD�U��z���7��n�Ǹ��#o[3����&��]���Qi�uP�ʴ;�԰��\��Ȉ�!ux���_%���J���I�uT��*���B��~����&/��`/	h@Les�h���T�<����f����@��nb#N�(��ஆ?_��/d�'+r��.�Ϸ(Q��l�9-KP�*�R�'��J��X9@�j+��ȇ6�qf��ͭeJN�c�	��L�I�����ҵT(�~����o���;�p��oRh�9bZ�ݜj�?ڞҟ%�ӻ�O��͖9�=�Z������vo��A^)Ȣ leњU�"�k�6����!��R�9I[RY���P���v�m:���͟�``4��L���i�;�al���a�ps4���?��H(�o^w�Nk�v�{D��'���ޠ��hb�s��7in��l��^Y����P�KK��e���B,B��� MԹ[��LK��17���OHj���y0������Gɞ��A7/�ZР�J�)j�#�9�cen�̻�k��g�I���xW� )���X�a�-��P���n�DK�u�J�҃�h���Ⱦc52��lX����zn�vq])�K��и�i��@ُ�S��E�	��r���ۊGP�F!<|�EPNI�!`2��*
�:1Q3�'�Pث�Oڏ]2m���LQ+̈́�
N��]�{�6���2��>d�d!X�7q�e~.7&G�u')�y.��(�Z�.���7��2�!�wXlxV64EB    1531     530�n&����9�\�D'	�������h?�$�]�N�2x:㗤��� ��e�KьE�����F��0Ξ'.��#Q�=/p��ꉩUw���o٥�����@�o6S�����WXx�}���.q�g�Hl����̰�U�+���KL� 7M���Qgh5/`Vu��6j��iY�u�.pV�����7e@�
AA�gQ��q1��<�粆�m��T��;�fD����z8P'3�c�<?�~)��3f���r�6���W��r��H��� (��Q�P��9�1-+hFe!�^��~�R���
�(S��[�!�B��p���� ��Ԓ�_¯�0}΀�5FGf$�gJ�E�����@j ���x]���4
.O�Ul�zʛ��O��,5�<oQ,�b�;��������[�/������􄍹�7��>��Ɓ��3�b&W^v��+�%u���Ҝ�26^�FV�E���`xwMG[������w�B%�~��#S2�f�**��Ľ��1�c����h�ʿ��OkĠj�3R����2�f̿T�-����|;W]x�����E����}�W��8S���fK��$��2Lo�����|��!����u���8:��gn�b����;G�|�4�>]{���yD� ����0�s]%�f}�b;��-=�d����'�$��:�$PN����h"���Y��X�֖:��Y�v"̫�i� 6��)�� �)��s��7�B���CS�܅�Ζ"؊ƫS��a7�#ú9�G�����|� ���&>�j墫'�5�����Glh樠���iF}���=q;�II�����P-�/O�8��f��c��I�pN;%���;�ɉ<j�������y"6:�~Ѭ[����]	�%x���ߓb�\�˃��	=�s%ar㋢��]�bt�e�}�&�3^�2�=�gZ�F��擰Z�>�xwd�؈/L���Dϯ;/����.���+Zu��9��:���u�%���x��TѼ2�]�OF��	lH�n�=U���3�@��>��B����x`��n��;ӳe��ՄN@��n|q���#˯�ti�J�~U�L>ɟWh-);�`�J ɶ]!���mjz��/kn��=Ԕ��<�8��㟣D[�&%0�w�R�N��V�M����p|�z�?%]���sc�ˌV0�]1Z�)�t-o����H�q�����թ��� 	���ߵw=���U�?A�Uӓ��R��Q3���Dr��<Y���ѕ	,"�4�MP��sQ�AX#Z��?�e���] �Ϧ����