XlxV64EB    55c4    13b0I�׋��FO5���eD=/@Y�m{�P;����=��<R�)%�1�en�jQ|J"t���S�<�d4��p�Ё�pJ��J���o�֓U_����KP�J�����{�c���n�`b�?f]6���$�_��/l�V�"���Ӎ*c�l��&c${&;iq�L���W
f��l��!�A���w�5�S[V��~��2���� p~��Ĭ�
�}�}T�mS����*s�r� f�mU�	G��2��j�;�ۙ|Ii⪾�_�������d#���9�#׎�~e:�a9��H�ڄ��si�Ȇ�����*�T�(����z_���u�nA�gL��.�3��g'芦�}7��,ju�dI������eA�o�K/׀��B�+�,^0�墑:�-e��wH$VS/9�'��%��<��L�~������d��\R��Sn���čݼ�t@�����B�r���f��e �23�ΫU]�Il���b��K\��Z؄�+�cw��[d� 9�{��A.ɫŝ�.}��}Xg@�iAt/����̏FN4����oq	�.�q�R&s)I�V��>�X��X�r#9 k@�.�&�|r#��Q5��8���7p3�s�%{7�X�Rb�;˷�-�zg��y5�e�K������0��0K<�����q�\���P��&r�/���H�w����~U>|�6C$�"���Ad�k��	��䴽^p�&@����$�ޘ0���yx��1�	�DxP\?��rY��p��Kg�䨲ز7�c���� a�0��緜Nzg��e7�Qp�����}�yz%C��g��^S*5��\e����|�R�#�SE�۟�W���x�R��-�p��ʳ��C/����6�r�aj�7��m}Am(�6;/�����֦,I*��»��mu��9�@JT������˾�:N�ϔ;W*�#q�\���ׄ���c���|6�u�G%/����Ed�(�\��c),��7���VJArCJ�y�K�3L�$%�iu+�BBFGx�P�$o�V}NV��p�u,�qt%O&>��<׵�0���L�,����A�'ڛ�S�O`���������]C?{��	6-X����7k�  �Y�*�=.���(a��fw&M�f�����*�[�~�(H=ԝ����ø�p�a����"��V9�$T�;�h�^�dBʲ�j�r���?I)H���jI��~^�?ph�F_tN��Z#���|� r�nN�Izw*�fZ�p���p�����#O�q�la��T�(���}R8�>�ť ��nq��i^W�������U����W��8f�[�áC���p�to���h��5�0��,dGB�U	��?��M�mN��P�qB��_A�8�U8��>�z�yE��e���hn&����=�7S�4u���Ϲ+�c~ۿ��D��Yn����ϻ�y�.ɳA$�(�?�]p>��vv2G=<H���������.5���T�*�!�Q�>��hg�s����� i��i1������=+�� ]m�_)M���0���I9�T;���DĜ���{�v��%Lj7;��)T�*L��8�Ľ#6%��PY��������Iq½v�^��-aV�:�������,�Uj����<���g��׫GR�^4w����t&�5.F�Y���H.�@JvU��>Aq:,ao�[a�ѶY�A�Is�ٺ�D�;J8���"�)F�H�<E�;w�dJ劑>���,�$)n�8%zb^��ȄI�7�r�k������ۣ6 $�����!�7;D�&����{��s��~�5\x�:���yޖ�~fSNF-wD��HG�'Da��P�V�o��OJ�6��f�p�u�}��:\��Tl]f/bA�v|�܄������>�xa͏ ��,p�4-b�ɸ)�HN�4��jk�<������ۛ���}&��Op�&j���(0����Nٽ &�K~�hg�;�ok�E:���ppG�@ub��Ço�_ĕ�W&k ���ڳ�����C�l�֛�BV[�?z��n��5#�f���guc�@�q�4��
I�Q�M�F�$5 ���s��1,��!���xH���20�'#�Rv��R�d�h�Ws�b=�b?���4!&YxoշJ��.4ʹ�A�������_�wR�d?zz��A^T�FK�$�t�4�v�g�F��(c���l�P2y��b�꿬eqc1&��Op|l{Ez!�/����Sr-m�,K�ZB���㰎�; �^FʴEY5[0WT:����"�DM����Q�z.LAF���scI�C�p�1j?����%O.x�[?_u�?\:��/�q����d?Ji�J\���O5�K�Y���R�c�`�:��is��-Qҝ�*D�$�o�~Wχ���ex7�7j!��X�u��l��i�i mW��d u�hL�,T,�1܎��'��阡s��͜5�g~+�����E�����W��`���9�c��Nr� �]��>K��^�R�$��a35�ݢ������|�>�o�O����$U�.��G�7"Z]�CF�����ƛф����O���~x+1.fO�6.]��6ٮ��T8��P" �LU��a��~�p�o�ɧG�_;���Va�R?�+�+1���~�3���R_\�t�	��b�"���צX��,�}����m��be���)��S�ˁ�5��e6ϱ���.b��A	+��H��'�q]z���� ���i<C	\�Ykx}�1�[>K�n�ܕ{��B��!����р�uk�*�Z1�����C��곲�����e�2V�x�;�͔D=XV���z�T`��j����M�0�����i�xbN$_�*������Vd��26`T��7΅bf�"t�	=�q,��x�H���	�t���OӼ\���Ϩ�pN���B�A4����m�'�|a�S�XC�b(q���/@�KyUM���^�U�}�w�و4@A6�Ɨ�!���œ���}J�(H��sl#k�s߇�>�C������0�6�TXr���'�nw �tE	kl�7�=|� ����}�o�C`k��f'0�+�m�1������tk�Y��J�fa[����a�[�.2G梤��4}����ZA�ڕi��|6>�* �&�2��9�1��\6��*n���%an��~�IVDͮ[x��,y�_w2�Y\~���"�r��rm<u�]�����|Ҏ/��	]?�.Z�����
(��?HY0��L%�e�j�DUg4R��5�9^+̫�I���G�ʌ�q~6n��`�v���X�Q�QY��y�Y9��U�0]�gw_˗���� 4��,Q{n�Mk�ս�?;��}}���z���]��K�T[�أڴ�e!0� ��m1:�qUS��l���?Ç�6�S�m�J� �A�!�@gn7j#��Rr	&�A�q�_��\7�JuZ���K���M׮΀�ʌ[
ÁKL���IZ�³�-]�4�vֵn�nw��
�+]�*o�x'��Ngc�F��HD���T�>%��� ��S ���!��V&E<g��ژX�65�Ue��_"�W6nag�{�	�fOD��"�����M�귩z!��h]궰~�q8aai����nĨ��5v7g��F[�A�QsLF��ew���ۥ�����	/.��fBݕ��L&=��+"�����o�/D�k�"g�V�@�c�g�!�l��H��z�V+�+q/\2\���]�ۆ���j��4�k�L�(����REJ�@��ސ?$L?��b����~X��X�4zO�:�L�>����_�{��Gnq�JZ�����w�l*��V	�x��8`��Zrk��̌�l�/����`�Y�iH���C�t��_P������Vxm�!���
�Ns(x��%��E����Xk�u�M�K���0PY��΅"�I�g�hHr�����hx��"�2�Y����1,����`\�,��A��x�I=���Li�%�z�$�,U��L[B)F�h������F��>J���O��@���,�#V�Y�җ�a0�꺝�G�A8�zx�3����B�PD(J=C͞@���� �C�Ǟ��-�+���}����o+!�#Z�I_QO9���0D���ü���3��}�;Τ�9��Ix�jH�3�d�`ёO����Gk{�k��i\*�/��� @v\�G[W����ō���Z�!I#6tG��O���~�R��,���N�"ܵ.7ڋ1�� 6��9�?�~�92��TطA��G������D|��Ɛ�'Έ����qΑ7�7Q����r��]�$]Sbc��ƒ��qGw뢫>b`[�2`�B,V�j6�<��x�F(�Ë��n!�\�?G�a��-Î�k���՛�r����=jd��E2�}|��!��
	B\�2k��m�9�`�o����s$��N��l��d�׸?/� �g����&z�AIV@�ZΕx�[���3I~-���|�+p��}�M��j��\7�R�̚�x"E�6&B�h��9�^�f5/
��<�/6(�A3�8�gv��q����Î�Ӥ�*Uϭ��t�r�{�t��Kv�~w��?�;�i\�©��5��y�|��a�?�Af�z+m��#�J�v�f!$)Gh��uc��F�FSz�I�������KtF[/>v�'�K`�|Ae�5�dG��Up�.@������z����Wq��]g�D������!&�H���G4#ie������-���9�(H�v$���"xv��g۴��/�lH�9�LN�H���R3����b����8}�OZq��&���!�1�_=���G㰳(=�)��>��\
�򽎔�r<�K%`%��c�b�v�S/'�y�=�����y�-9�7�6���m[����N��ױ)�j}��N����������y�+��XH�x������#��8�6�߯(1HɈ6_��_��I�;