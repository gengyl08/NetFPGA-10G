XlxV64EB    2279     b00HcxF �]\5Bm)���h_{T<;I>8���`�+��.���|�+N̗܂�����_��]������zT��xK���T��v]:���%��\Q(;[����=��`QQW��
�T�E	�B\�� 1I�E�yC�x��(�t��f�1�F�þ����"�r�
�bY�L�D�oci�F��'���h���3o%�[K|�w����
{~T����WFoWԸW��R�L��(cU��m�34B�!�4h��[n@�L7PƘ��x�C�M�����T����t�͏�\��:�����,f#�H���^�[����A -�aCs��C�:�6?w�E���:��<}[Bvk�h[l^U,*o��PL�z8��+��0^�Aж���T��!�h�50B�h���)%7�٫�����~���]���{Q�u��B������gS(3v��{5�,�Е?s��/FI��p�@���'����Li�?S�H� _g�z��S�@첲C�_�/�Lr�uI��T��� L<�HEP������7�����v����O�{wdu&��̍�P�s���ag��+�j��p���
oA3��{�j�#O;d`qUYak3'z��r��#����3YAnqffQZ+�B�C��?w
����PJ�ly�r;�w���ʼ^����A�/��|�jv�m����q�0A��@��`���6C�������V<W64�DD��J�)����S��E����Lý�S�[�vutAB���+	�$'6B�֒��.=�2���꺑��9P�8}���TY^�Q�I�H7f+�/�cAб#�k޾��C�8N��&�&>���Q�<��앾��g���Wy,U���pO*�����I�κ5
�K!$���9��;0��"Q�=�ݔ*nNl���*��?��]R9��&�NфF-����)|��"�Y�
�	+�p��������r1��#P� ~�I�=<g/͋��#%�6��� ��FR��Q�-x�~��W �D��0a��Z�LG3Fe �W�ő��J2��3��Fg�ۃY���($��PAt*�]�8]O�K���ͱ@>Ap�'��**�gsݔ<mfE��
�6���y��G�Ty���'��]�sT� �f��~�`|6)��DίG+B1Iv�P=��t�����n�"!�W�/`��-R�j*�Hha�N�ą\e�i٧-�P%E���S���B��?�V��$�v7��Ltשl� ~�Q�\�EC��u�ꧢCMY�U���S��X��̛bW���ίπεQ}�
P����{^NF+���6��>��y�ޒ�b��1AEW�*˕��4�H�_uǓ�lG�����NQ@�=�y���K�~�qv}�O�<��XP�|��._r�{qRDu��,�v��o I��f����d�a���P<Ly��,H�'_�Ez+.߁3�@; ׅ��� �F)�k.wǷ����:͠ ���A�{h�67\ՠ<����Sm���a�O4�lhs�Zq�}Gپ;�|��">�<)���V�
*�u*w!@��\D�uGV3�X�-����������9��~�(��k��� [jJW��Ov�1�����ê:Nc�EX�//�WO��d6���qa�n8sͽ�Ԟ����P�cK�����w_RP}t�_�UV9CDS���Z� ��h��J*-_�S4*�~O��=�A�����
){��.��3,(d# ����L�Rɴ�4�����"�yl�ɑk���zZ�T����FG��g(��
�	Ӵ�:վ�rxr��Y2�%#�:�/t���q���9nV{�=���q���+k:̧R�|<ȉ?�bJ6X�m��`�
�� � �կ_�^C �b��^�v�A�vw�}^�����_p��,�2�$s�;5�ʒ7,=�6s� ��ʔ�,Ź���ʵn�XN�{��������a3gB��j��h�S�w+�:�?���gR5�-�]���f�!��a���<n9i�!:7�|v���x�A|Ҳ<;�!��[�9��-�5C\�E�i�5�HGk>L�[`+�h��Ю�rq{ԁ�!�YW���)o2�@������0C,�]V��G��6����F�,����nwH)eE����~n?�:����.y@=-V7�j�^I"���;�K����V�s�Ϛ�X�d��Xt���81y��a�sI�yeْ]k���`FW���ñL�ԺRp���L��\=�OpW��46��^��4�����cV�ܴ��hg�ʝ�F�w��m~�[���H(����^�m�V�-�}�3�0|9!�+�7�*�
�O.b7m��F��UK��ն\�y�;�g_�iИ�)���݌�t�*US�9'���\ߡ%ۅ��.��>b>�Gnu���3�R/���5�v���0��S��38vs<t&h;1ɗ
�T5έ�r�H0`�3�+hx��o;C�&�#Z9��N�]��m\*[��!���e�mh}t ~���@!�]�Y�da�!�<+�'&X�O�B��l�`L�|H�Ajl
c�M���;]���X��V4|�` SP�ȯ���Nu)�\`D5�b�@a0�x�B�vZ-�
w�ّ�e��r:�l�O9���[�%�v�2V��@s�%�@���s�����8>��պ��G[���N)����%��x���&�q�筋�����ȵ?�m�yP@���{4�M�:���k7���$x<�6����-X����ָ�V��+ ������m;N�����ȕ���1��Cտ/��Y�σ����MSS;��}�Gv���Q1@Cf�#/�|�iq}}��x���