XlxV64EB    191e     9b0$��˽�ʇ���m�mu{��R�$5S�kY#ݯ�_�qϯwȫ��ejCq����]1�&<�`=��u�历~�ӴP�~�n]z���F��8������J2*�7���G;�k&��{m�e�c-�N?�Ǯe�5��y��<�mc�#G���=��Ln�05����;͙L���9B4�pG��S[�M����KM{�P ReV�i5ct���Vi�"�&6�H���r�d�Y#r�͞���E#D�������QK�g�)_CE��kz�=
bU�-*�&Y��7���ހ���x9y��F��%b_S<Rw�6�inp/�L�C\@\��݊�Ĉݍ���zK�]����Y�o�3vl�\��"F���-��6y�	�W#�j��ں���l��_�4c��p��&䶽�,F)ݚ߷���)�_�ڲ�@���|3��1�94�b*3�%�+1iBb��ns��:�O�{(����2O�"!�l�(R�s�
�ȅ���N������!T?��L���^	(��A7{U1�����k�5��2^f%[��f�ba�p��늁��±�(|F8�w%�G�OQV*Am�}���(IP!��!����#�.�psC�
��������uFG��M�F����ch1�@\sr�.uTq����`���E��Z-�N�R����Xe�
����1+:<���f�� ���lr������ڹII�:�h��5�2�MLՆ&ͨ��W�S�t�C�8�0���Q|۔1k���B�h��9�
����(�D���K�Vճ�8��h=������e ����`�[ts�|��}�C)�/�����W�7�I�=��1��7�,��m7";�w��·|�eN�����2����.#镆o�'.�K�����T?ѫ��;��4_T�$r������f!����̚����֨5.�ԁP
�A�"h�Β��P> �DG��54�c�9��Y�6��RҶ�ϩ�=�T Fo5�zbӓ(d�g�t�hٔ+"��A�L�	<�盵�]���Ti�'�bSЌ��
��4�� ]|��]Ҙm7wӛ�W��Oqg
�Dc܄��i, �����Rv&z���Ș$/��� JV
�~��6eƢ@0r��I\����q��4�&l�[3�����ù���!� ���ѳ���s�dH�6?����c��^�EJ  �	�D��<`�N�Ci$<��v����a�߶>�Ӣǧ.�6�/N)�BЛ�3n�M�SO��q,��|��"(F*^����~�h����6����ݐ�x�����lw���̰�DLзdT��\z�ËX���S"'P��"l�y��rhTXi<�f_��9����i�l�~q��(�&t/O�q���m��IS�s�mY�}���}�a�UsA��3������)A�tBt��zdDi9^.�ۺ:�6���K�a���( t���~#8,�Y/=���&�v�I6,M�#@櫧���1֘S�W[9�����X��@�1��|f�)�!�b����2��7&�WI"^��}��,Ȣ��ŋ"��tQF�Ӹ�������ѫ�KrRT�q�'��N���|�<�H�JL%c7�Rv�߳Qa��'~%U��r�Q�6ٟ�����Ք��� ؏�}��͉FN>���J�c�a	�i�eyQ��$�|����� ](6��ԓU��Bd�}�K(lw���WJ��_H$YG��RKȖ���-��3۬[I;���&��M?X�EYb���7#:�>8��G$�
�~���!�b�mG�� TM�?����n���9gR�����W{��Q|�A"��
Z������)M��F)�[�j�ն�~,����a��'�X9)�-q'%�����|���K0�4�X�1�h��U�^2V����3�^��[�i~6�.GQe�W��.�E�[�)�
���p�2tVS��O����;��@�}/�繌����Y�?��0h9l�b�n���Up(ƪz?�[�/Ӽv��I�j��/yY�)�V;�N�P�o�&�%Kx\�xΈV���	�\*}�x��XwK�~+����F��VKA�z��e|�,������БC��F��xqqA%�X*���b���V�b�C�S�RyC�M�J_!L���9N���]14�6�J*` 
8&"w�ӳ��,㙷�7Q�K��{�v�	j#�I��@X��D����J�>_��h�k
Q�=��݌��`���EI��1"�l�͵�����j��#�%��Zr��αBU��S�<����k�Lׂ&^��h�w0O�4_���������YO5�G�TR$'"e !Iw���1�����?����B��V�#H�W�<�g�'5�iB�pHU�栂3�����MJ�KJ���-jm��w��&��-��_Η���\q,�3��������jF�Y��:�Bn��մ1�Yq���H]�/���-c���I
�mCY�a��A�>���rJLM����