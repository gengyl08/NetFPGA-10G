XlxV64EB    4831    10d0����!�V7X�_
[�)wp��
�q�M��H��ٔQ���R�4V���	~�^�z�D���sh�b��s2"Yqoʁ��Cݓr�}yWq�`a'=om�//�XqW"�ɻ��B����9�AS�s
�\�ӝ��ќt���u]Qd��C�Y����f�^�뺷H�'�ȑ��2i`Y�@��u��A����ĸnÁ��\�t��و��=�bzI���&5�*����omeg��r&P�ǻ[ɓ�Ĭ�i,��^��LT���sm����2����٬��^��Q�]�qu�j���z)�O�,���x�2^�Q�OmZ�v����1jl�۬�$SMU�YA*�
���O=F��ƽأs���?w�xn��N��[���ʃ���Nm(*��@d�>���ξ�j�#�bi�E�r�.���g��X����|�Q-3N�0��ks��h1�܄����e�`��#)���,�-jY���@=��� �B�/Z�r�^�������W���d��R���#�B�K�um�4)x���⸕���N�i-JXH��@(���- ��:����}0�O�4~���$��܈m���cDr�:��'��JM����r�d���bܪ*�K����@�{T|	��ߩ>�?u�׼")�Yt���O<�.�j��4�ؼ�s�h-�r�<���}M���b=�j�r��7�&�ţ�D��丆O5�C'�K�W�ͮ�A���-�g���i�}��ۿ��q�I,0ek�	�q˸LW��xETlBO�������8
���@-��U7.<+��R��w3��*���)>ٖ�lg��z�u��q�R�s=�b3�J~��@	��sX<�8�:L�'8��+�����fP�'�_e�۟�fN���!�r>b�h��(`�
�Y4���-�m�����ͽ9_I����>юڔј��O%W$xZ�ŪU�"*�ǒ+���;��4����O�Q<l�HHW'�IS���	W��+� �uDfD�O=�竽����5�1q����Q�ű����mϷ�ʆ�ϥ�����s��Ӽ�?�&�!��."V{+$`<�8�n�u�`J.��O��L懕&<qt��d\�f�(N���#�!�4'���=��7�)@��V��=WO�h���}�0���?ڏ@���E���q�YG�}~q���0�G.8X��K��i�cLr�d��N)DDYO4�mN���}�4O��=	@Z�T���D:1�����e�PW�sך���`^����G0��4IL����ֵU�Tvԕ�����ĉ�>��Bz^pԄm-��힦rȃ���L}��걷{>� ڇE����e�@:9���S3j�څ���Hj�����w ��|���XX48S���� ���~�a�n�r֯�@��t�e�cMj����ْ=VC�l%���P���9��с�Y��������hqE#:�P=�q)6�+�^�k���ͯ}��i���'�ͯ�<��[+���H+�ߢ��&?��U�1)�KUswBCKp�������v�?,kJ6R��.���P���Q7��0I|7�pL�t�8��Ї���5I@?���qoy��W��@��㎾���*g'y?�w�&���ע�6�d�X����u�1��� V�C��ʳyW�:�/��rE��z���s��t0���Þ��ʟ*�� ���ǥ.��:H���n�����+h�	�]O3qj�̻�z��E/a�bW�^���W�O4�b���*(d�K�O�������[,��k/���ݬ�I�=5��F 9%�V\�+G7(��o#�b�=z�	�����6M���Լ�	�/���ܯ~A��?j��9*��Jy~���X�_��������e 7j.��΄&{���:RT%�ރ�}����ZX���I9aX��5��	[�,h'�4��IkE�%~�JƪY�A����k�����ٯ�]�h��2·�Ћ�9&�rMRN	_��w�ʀop�O��@R�=u����U��� K�@?B����:�=�]鉊(b���ʘ@rg�)�	ri�!1!RpN�5䬁˻x9�`U�h�"8��Sex���q(⬙�=ꭧ�ҭ�%��_�D6�ȱC�2���#�6�i��W��m�h�ϞF=l����f������қ;�*�i�kE�r$L%%2�Ә�6�uT*�&�5;��۝wy���[h����n��Q��%�M�0�C�t9��qP�	�ѲO)g����t���K�W(L��˳��G�eb��^�;��!^QO��,"���@��肏�Wu�-~SKI�8�j�v��/���N&�z��uڗno�h���T�IqN#H����H�!��ht��1W8�ُ��هZH�\םRᙽI5ֱ|8٭�w .6FXNx��3A��nɌ���Ǡ���Fu�?����S��9���N� 9�$��v�~�?G���Λt����h���<P��+ B~=�V�g��ȟ���q��*BmV���)���y����ߧJ"�ݼ�]�*Z��k-��a\�a�s�P�CCOӸ�L�"U�^ ��l{�{Ck��-W:�K�aے��>��ZT����&s��H-)	��'2�F�M�h�}ҡ/Q��j�l�v��g� �즍d=�Ҿ�����ʴ{X�+��Yzh �,X6i���u���t�M���T,�{2^��?,��8e��6%�D��&�^ф�XQ^"� ��E��1���>�߉P+J�cT׎����Y�� E�@��Tz1a)ХeRmo��g�\b��jmR�2&i�/j�>�2�Iu#�ύ�ur�5��|�A�3_ΪiG��$V��2-A2e�D�8����l� d�$��5g�08y�]��Դ9�B'y�3����'��]����Y�!e`&G���!y�ӰT�l���T7$�8�+�rh�ն�l�&%� �	� ��c!���Ⱥ?u�J��*%�C��'ӛ�Dn�&��Cr`Al7��yȷ��T�����?mM����*r Nn�iE��݇�xh���5(L��|u����߶�B�l[ȦV��@���Z����B_�y�(q�"�9]mX>�G�=J�5����̈́�^(�t�:��|Z��b&]�BO}����`�Q�64��`c�r�q���<��?З�)�1�1�G�i�?�$�nm�8ݐW��8{�����v��uGO�����|YqC��,@�1�,D�L����<���fgj��$�.���SV�=���rl��qѕ���q�󅙆o�iG�� d!xa;��lϘ�v�d�*J��QTq}�X6V��}���Ѵ����"̚K�{K���!ފ�tb�z��Xd��y��Ƃ��ڐ%��V��ֈ�?�
-"#'�$�L�q��=�H����Ȝ�X)��돁�h��B��֖+\]gC��S��Q�& �.��I��bY�y���!�k���6���f1?"��KW�,5��'���4k�h��	lǫ�#Sp��m��g���MM}�_b��4�k0�,�Uv�wC[٫Jj�O��A�u��G+��2� =�*	����;Z��OY�{��r7׆\�x�`�ʶ��y�L��N=��8srw��u0D
�#���^���Yf��&�iu��w������m��>3��uNp����R����"� Pv`N�:�!�-%��x�3!E�J��0c�UP2d}��2�h�R���(��$��(8��2�l�=�~^ѧ3�Ks]�y�ev�k֑��&���5!�B�3�u��I����.�����{W��+� ��U��(�
v�ݺ|�ҭǖ�m��O�,�|:�T�q�̽Iy�>a	8kE鴇&	�$6/�]���4Sk# �����F6=��&k�M3߆vl�B$4�o�F˰���%�,S������ V����� (#:I[2K�:�%���&�0��
�Л�q��F@-
=�*����d���u��l�UK����m��q��V�3�wgm�����T.���Y`��/3zJ8 D��P28��&`K5]F|쪕�(k-��ʑ�Б� ��7i�A���jn�?���U�Uy�l�I��;����j���L|cg�G����S(P�p��k����:+���v2�?^�x^�p��(�����!����_���T��Nʂ҈Õ��Ya}�S�ߒ;��	lH��0>.��
K �q�G�+�*h�{|�{n7J���dX�l3�֔�%q����V�������W�]i��\�N�t#���U�
���0f�~���>���!���<�$�r�����h�\�c&�c`���2~�v�v|Y