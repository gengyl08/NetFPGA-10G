XlxV64EB    1fd3     ae0�,Nƅŗ^�I�̙�I�9�i,��<�
���ۍb�2�.����2����,�pr�nnt��&s��;¦����O���!L�ַ{Vz0V�)��,{���J��Y����T"R`���Jv\7����v���Ka+߯sU\T�g|Y"L�!ΩX���������Yxg���>��	6؜�����{�[�|u=�Qy��@Vu� ÷��8enK��/��y�6��X!�2��L���б��,�X�
\(���>T����o�W����7�kȲ���{�[�1�fk�FK�[W]&`X*̞z�T���j'��'Y��vҡ�M48�xZ��Η/�F�~r�gIJv��M|�u-���_�B��h)�y�j�J�XмG�|9������f�{�A����4�N�H<S^��7�$`��$��>�#*�,�?Hˀ<96�o�ef����,* شN�l]����р*����N��/�oh�`���C nv���Ϧm��E�N�汨qht��8s�3[��w�Y���K�!�k��ia��_�մ������|2�y�ц�����;$´!ۭT�GlLޝ���.,�|=ˡ��)ǻq~����@yV8w�l�*_�c'���
�S>��pΊ��]i��/�S��3Z�L�0��l-��e�5=��3�r�M�k.T!��.N]�w��J	���j=���y	��?�\��t�T{b�LU��
=U�{E7.ϠR|�7h]�����S�/�מ6}�h����=w�S��C���ޟ�a�[N�1�]7pop{�tl�-G����0��Ț�(G�����|Mٺ9�Q�}��� n����ֿ����{]�ц�7����I�Ҫ�j!Z���d$����T��,�-	�o��U;�gӝau���*[�fUn7�B8�f9TΈS/'@��p���g�:�b\t.�(��W�K!���������{R# ��2+��@2�qMS�Dp�p�CT�-��e�� N7��w%�G\}�"S��N+oj$k��'�7����A��YǛ��o<���Dh���'���cĂ�v1�4���w�t�S+6��fv�&�"H!'��W����U�u�O!*F��
�[�"ɦ�?D�3�����7|+C�'�=��k#��a"C�)T�^~��K�;�\�Gw����ծ�kC\͒��[j�AoW�"�4���{�����3�4 8A�,Vb�XQO�[Ɓ/�9f�W[V<Z�^R=�G���+�;����e��8O���m�ߌ����<�K�;�F�f��2�۲��P^�`s]T�X�Yמ�(�lҠ<��e�J�d� U(j����C�C:�s�1���]7�^Cs�7��;$l�����\;g`�K3$G�ڔ����Ac����� ��+|�]�k�'��q�ܼI5x �ż��F?v�.HO�˴L�a*<��/� ����.��ܤ��`&{��:;$Xt�u�� �KO���qS���Hu�k�c?wq��گ�`��w���e?��
����D1^y3�@Zc��B��$�ݧoQ&��\g�Rr��<)�N�����~�%P+%{ro�zVN"��B�*���6�V_��U�iȡ)G�M�A���� �g��[��UjN Q#Z�8c�A�Ј���������$�m�(���o�}�8���ꑑ=9��ѦI�"�Y���\n��٭��N��P�6̤ch	�n�2�um"�*�sh�SWU�L�\����pΎ���_%���߉/��A[}� ���ʀ�K�]�.{��m��JT{OD{��f�^���B�~y5�����u��<�Zz�Ky���_�L����Xg!'ÿ�ՋT���0�@��(��J�� ��o)�~�Zs#�I�W[�s��r�H_��c����m;I ����3`5$����B��-S��%x���g����5�F�.<��B���BF�wLu��0k�-�y�%xs/֊_W� �d{��2��`%��O��Lt9���z�q�3����`Ѕ�/�u�����VM��o��^i%�^��@�����5��k��X`"#`^�Y�f	�=gҹ�v0Ms1iá�� lg���9�Wޮ\��j�O�ð���h���R�c$��IX��$݂�6��Wpn��S��π	y���ܘ>`1�������M��.b��,��\f������]$l��B�*�8K!�(�����I����ֹ�`c��Nh��@ө_�j����fŦ�媁�Dȡ��k�7k'����W���i�+K-e��qD����cQ����a�M����k<�����(Uz[��n=f�h׸���.qE�m=]8j�^�{L�.;�VF;%Jڳ䱑�tX��R�"��,�-��-��2c�?ܶ^Zx���6���5���,�򙆒8�Fa�/���{L�r��$ڵ�Q�f�MU���f����i�Z��X�E/ƙ��EQW4�Y�p��Z7H�i������u��J������أ�G:c!]�F�H*|�KP�ng@�w= �۰D�}��h~��x�rX��rwa2��~$���w�[��PF�
⦾�ᩯ��S��06,��Ym|���!>W�T��;[��ɹ�_��б{!��)���3�^l�w�6����/#'?���f.m���f.<+�c�+ʏ�`ي���4���n�o��@��0���>���kx�@�~�D#�n�q�15l?�t΁�R\(!>[�����%�h�