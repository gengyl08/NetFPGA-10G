XlxV64EB    46a1    13d0t��4%!
W���j�֚˲�'��~��DҢ5�A�h��3����UB.~[�W.�Pf2���U�z̟NE�1Ew�E��;\͚D�Z{�C�� �r��@��A��ʧf��p��=�ϞD%=fYczϐ��� s-���I9p�Mµa���Ŗ\͙�,3q=p���Zh���MOjgF�H���~�G]�Z.1x�D�nD�}�6=���TY����G�>�;�	pv��x���V7j[�i��,q�E,
&�Ď��X�\��U�¸���������<l�	�9�ƥ�fڠ����"����cv��[��m�w)�,!p�E�d�Ɂ�������,m:"��f������������M$�����8���{M�k��#]@���(�`Fwrl{2Utj/�`��ib�D'���H��x����>+�{�muwo[���GH2���oobl��fL�3 �EQ�Y{����#k�׹xxI�2iu�c=��ܥ�
�?כ����<M�v{��Sz�t��}�Y�O��l(�2��R�(���7�&/�Y�lԕ�B�;�&�c��x�	�E�v6(f��jx�0� 5_�w����O�)�Ү�'����hT'������[rUܖKP�
��@S3�l�����6@Ǹ؞�5�'��|�ሩ2G@�qQ3��d�QX��$[��wL�?3@$�[`�	aZ���{rB���5d�mD���fE��3Tt󛩂�f�����)pZu<N�'�PU�sy� ����F(����
�.یK��D�;Y��]n�Y��!HЬ*e�/"O;�3X�K4��\()��W<�s4ё>V��_Ɠe�k#���8���_���ֽL���af���b�i�v���o���P�Ν�E��N�e�A��2�H�1��P[\��T��PU�,o�\���W�8�w�ԥǑ��9�z4R�X��	�$�j��5ꦑ�̖�I�@�p����$h�R�2�;��|���<H	`�{���v���#zT�\lU	|c�Bk����i�#�f��'���e{��^ϯ�f�!2c���t_�r��a�<�Ix&�:F���7D?m����_���^AM3fr�����K<�C8��߿�!���N��bJg��C�&a�RW�#�R��GF�q �/,@�ùZ�\�~ѫ��W"n�C��x-��{�̏ε��[0��N턔��-�	/�ų>"�2�xK�b��9��S��NidJ�0JR��u9�Rp����rܰ���I_��4�u�ڗ~�_���݇�a���QF���!�G��?[�i!���i�;Q�� �Ā�d$�S�a_��a�o�H�;{Fpl����,-�T		��u�M��=��O�1$���%a��;V b�o�!��t�Әr��qP�P��eu:Ȫ=6�dQ���S�}�V;�Rϯ��#�_�@����I�Q"�2P���Y��y��0���YFk._�;�_)�u��?���^ A��n)���eQ�q��K��n� �՘��Sv��� m��G�8�i��õ�1/U�a���
U(������\���1c6�*�;p�B��C����
~�����!]�����,]�
pg0A�Ϥo�8�vq�A)���51��68=6&���>h��-n�����#(��s[K�m�0t��"�3�}l�n��E�$Oq�?���-�<ˇ�����y����U!�yc��q��ݐ�`%?��fe
��J��z_�4 ��
�-�_[?�4�$2�}��b��F;	<���H�F-�O*���:U�NC�N�6L����Ղ|��Bn�z��8��ۙ�ƹ����9�������[+���}z�(����r����`����PTKuq!҆�r��N*<q�B�/az�I*���f��b����>f\�kw����caH��]�T�pZg* өB�h9�z'"$�4n�zt mb��F��忭�u�|��|�qFv?��l���H��a�X<|�;�����[��, 1���.[L�� ��h��c����Y(ٛ-�}����W�d{�{2�&˰�?�P;8�a����xD�o!��Ъ�4����g����PR�T��0�wp�L%(@���#̝0m���%���r�r���#jJ��i�j���C5I6dl�3�}S����"����L�@(�*���
6��0�p�z�\�6$쒎�'���d��+�����뀓���v�I���=-@�fE�ޗʱ�R�&D[��xH�RN�Unr�������y �\�A.v	~ɗ���_��p��ّ� 8�b�9.`��e���� ����;�����5>�����r8w>�۶��˫��΍�1.ft�&�ֲ~͢�I)$���b��D���w�z&8Y7�$[��{ �WN'�ӛQ(_239���������� ��H�'���};\����R��"|F9�w�u���V�J��B�F��q@9O��o��\E�	6�a}�0�7h�'�@úS�|�*�9(��W;�@����m���T��S��
Ӄ��
���	����밳�[�ܙQfK�N��YY���Y�`���Ϫ)�����Z�
�{<q�a��hr�Ы�-�PQc�\�����b�f�0��|�4񓦈�̾/F)#IC���@[E%kJ}s���Ya?�l�;v]�`�ӫ���y�E]`��������?�F���\��9b��!w�RFk5����j�Ap��`��Xt�!��r�XwM����`�=�Mٍ��J�)P����l��@5�^4k\\U�zC��c.�e��d�ZϦ��&�9�
��'��ߵ�J�����']Q�h��1�Ϗna&�P�~9=����jmߨ��RC#VM���8#��H�����(��LpF�=@ϳ�����o2I�m�O3G�8��C���Oc'JJ���73�,mw=���U�1�B�F�C�g6I�{n} �$��c ��I����I�[������^6����WP�L�p@� ���h�ԕ KrIZ
����2��l�CK�WJ�K�w-;�6���Z�nH��e��퀄c���e-[�({9#o"��!kr���,w�LC
����E�Λ���f�_��S��NGv\�'O0b\���r�],E�bƬ�H���3�˙�e��?b�/�-
A���Ç��m{�7��e�B�<;�ݎH@/�QI+�p���F�
r�xP������Q �L��vi�b�DB.�ȡ����0\,=�e�=��ǎD#��]Q	��ptEC��U��պ�����y��ŋ����
} ����Wr�D��D�oQ���)��8t��R<���S���i��ce��?���̗��R�j�t j�kZU\�C|X 9��N,ڹzS`!Ζ8WtӴ`�[MWmI�B��p٧�`��
�~FUϧ�f��t�Ŵ
F=��t��F�r't=��0�7CĪ�_�=��^Q��V�N��6C)Y���&P�Ӂ�M��ɱ�A�������P9���̊H�5��o�ނS��f�VS���8D�]o��K��]_�����D��։<���{���,\�t�A�	�wg��$���WƤ;_�X�5pwz��H\���I��9%��0⍓
.��BO� �b}_�#��f{5�%��~�'����q�N>q�B4	�{�e"GFL��������(((�ۻ�la�u֢_j}7��dʫ�5�`�ع.+ ���Gu"�d-ݹ��7�C�[s���1����>�ޤ���>����4ǿ�i�4�.���iC^���Ǻ(����N\O����X��1�z�p����A��Q�Q9B�݋Hר��P(�ч�+叕�b��]�|��^�5�ߵ���I�6�َs6Xk+$p���Fy�j��*x�ћ�Gy�=��\!�K,�ad��KW$-'a�)Y�^��
�b-b��Znr@n�t����S4mN�����D�Hա52ްS*�!�yM�� ���DP҇���˓���;���r&6d8�X!���:kn~�����ڷj��$���t�F�0/�r �{m�)�%'�VGFe�&�hǌ3?U�$���@���IÏ�_R�k��3�x92�NX�^.�������������Ӵm]���̞�s�"b��:�ǣ|�ؓ����Aẽ-M6�)�D��HY��Dy��:n�hs�P�e{��bb�8礙�9�.B�r��p-�������(2��S�3,������xS�{��p�G�
��\��fM�\v�&4�_wF�} �M�J��t�.��A����@=aA���s���M�.8�[�#D������͍P�W�2e�W��]g���5!��d��I$����%�ԅ�|��d�u-D�y���Sy��`�6���*�ء�NY ��c��4��`p
��M�#���0Bc�v�����uH���S<�n���A;�c1��D��.������i8A������A��dE����:Q�������X�<����J/`�h}i��٣�$)���#��F} `�� �亷P�*)VSfo`�V�w�`^�\�Kr��w�h{$zD����T�/�ñS�/jUe�Jͻ�~�񳚕��i���aO��tDǰ��H�����4�'ð��':��v�3��� ���}t1U�l�H�-e��]sZt$�����i�M����46�o����~k�Y�[�[���5���cv5�{��G%�.���:	둁�b_��\��CHBlҢ�~p��E��ՉG?W��$�Z�"	%��%���>��˂[T?:�E��P7M<��c.�N����e6��m��ce�r�Ҧ)����1'�6{����B�!X�vX�o�Fs�I�һ~|��������o�����8n6�W!��g��qʝ�k��IB9BXƱ���Q�9�({�pb���͋�"Jƿ�m�����-�bw�!��-'�O���g�+���1S#E<�����9ղӤ�~�G��=R�^���~vg��yP5Щ�F�����ĸw����#	eT�xB