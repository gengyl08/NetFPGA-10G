XlxV64EB    3361     cf0�59�>���5��r�O�:Y����@��0���<��m�/\n�EQ�ê���#���0���~��96���,;�V�I����$��ѿ�`rb�{mh8�R@��H{�8���^C�,r�4���"�e���V�J��A�4A|X��2������5m#�d<��OOA0z	(�2.B��΂�'��>�Fn�W
�2�����m�I��C�/��4��ħC��.�8h��u�ʺ��GHd����Ud��-�ᚄBN�d������Z����钻��F�'���Y8��"�.NZ3�7�z�t�m+�]0z���3q3E���W�q������MZ���p(y�M��z">`8�����s����,.c�dJ�T|��w�x������i&���k���	�\��M���\V�Xh�Z��<��q�=��8��-;�c7"�,B�Cj�v�o���S��#/��S�݋Tza�r�Aۆ^	���u:ZUN���q�>=�Po��o�ʲ<TD�/�Ӈ�΄/�t*�(��"K�:��qp�i�hn�_ 7�-3�C�$%�^]��%I��'-�G:̭&��]��\��T��E�
=G�k��r��pf���iu�В�O�KEYy�n�?|-"�@�'b	��A܂)�zD�G�����.��n�v4�Ol{s�b��EK
�.8���D]�Rv;��	����,C&��"mV�VzSԊ��6���P���}�J��I\ĳ�ƒ;�hIV"�fs��\֜��'<cW�,�q:����H:Q����a�0a���A������e�M*bOߟ �F�]BI!�t��g]g�6�O��
�K�԰K�a���V� ������հ��
yJ�Ş��K����ŗa���ff*o���[�N�EG_Џ�����9y���a�Z��Z��nO[���������hk9U|Cq��OQ2���pzn<�G�=�@�`��҇�/A{�7rr�T��B�ktX# 9��R$�c�>���};�('���(�@�8��G�<	��;6~���Wϭ��W����T��s��Sq����-H��;�L>v�#�1e{�9��P��||���c�u��5em����5rTpG�҈%�����|��<hQ�/��O���{B;J�>mv
᬴�E�;v�@�y�L��(3��9)�M���g�ciAL�S͊3��0�ͮ�����Pk�|�������
O�)���x寮�)�~�q�c��1Nnv/|&��I`�"�Rk,��;	PE�Կ'�La�K��aY��*��W�u�^�x�w��LC"$��0Yy5ÅL�+�7�gՐNTT��l4�Fc;��̔.n�Hc	�Q�O�e��D�$t��5����#M��ȗ��f��h�g�oי[v]%\�)h} Z�C��Q]�a�`C�_u��L�
�
v
B�H�ca��d���j���x��Xd�x	)��JL�/�#�J_�^�6m�
fK����1��N��E��,�9�t�|���*��4}�.+-U8�9�rx.�'BK����������}�!�����'ݔ6�P�9�aNX�Q`h�
��i� ��M���M���X1GDp�-s$<���׊��G��n��YJ�µ�K�fMr�"J��E �0��V�i�7���Y��~]X��|w��S����+ %f�		�^8���p���Qz����TN���Qפ��=���p��-W��yOVH�0mL�O�{ ,a٬�M<-�VA"��ƫ%��V�&��R/"J��쫩���&�c5�]Թt �=�W�p��E���<hU���nu��@{k�ZE���l}o�p���}�螰���L��"\�<�5s�b�D������c:%4e��t�W�J���i�G�2W�"K��Rΐ�B+�hխ=�?ļ? R�"�C=R�}_�6%_��o˯��prU�>���vh�-Gӗ�U���s�։�*�5Wfi��eOSc�
@i{�(.��Ă�@��ٗ��c�^t��t�g��O�i��#�d���?�O�2{O�:�2�@g��!��n'ڃ��,���O��GD!��c�u�`٬��a���T')�KB1���B3�v�	R>"<U1�\�句u���F_���C�u_��<��"��v���z�P�B�p��G�9��	��W�kN��(�&Yuc X)+ ������#p��=�D�%>���촙,��G�#	k�&U��s
�^�dR2�Ά�(��VX���p�W�x�M�1pY�ͅ���E��t2�j�FmN��6l�/�W�-ϩ��e�Y���l��,�J5��Á���Xn��gg�γ(�i|�P��kcc-O���������jԐ!�C����8�1X�Ԉ�),+��v߆�7\@�[�)��6/y�����Ss/
@�*l��M�VV��Ib����u�P��G\��ƋeTNW��* �����a�$7i{���6�dΪI����à}�W�7}>1w�"d�ݵ�j��Ѧt���.�q�jz��ws��g���]�2��݇!D\����%��T�s/�ц�+&G�to��T�	�_fI��h"O�T�޷a%-��@�8�FJ\;�h�J��w�h�u;���2�q-���,��sK|ESb��X�8f���D��3���As����)�ֿ�����i\˨���2Ԁ/@��Gr}�{�:�P��Kf΁-"�_X�"�޿���S�����;�gy��������L��s���ȟ]){!��W�!_;n��fl(�1 �4��Z�$�.��:��U��	ѻ��������H��ԟ8/c��U2�9VW��{��Q�+6mAe�A�����p��� `��V(�VX�0�`�	&�9ÿ1t�\��%C��K�1��g�c=���<�˨�.2���$�x�9�������%~�Җ�x���}B�Y�������0+>'�'���7-�/iw����Y�K��]��7��0`�HrR�@���	��Cgry���m6J���?/0��ℤ����ye��keZo��,[�a��� ���5q��ZhF��䐊�F
��A�;w����55�;=��/5_�n���r�F���+��D����[0٥�X���� ��
l�(3s��TXX����B�P3��^�
'�V} ����7v�FHcnc[o����`ɂ��2��O^
(p��M�-����~ �t���[/���hA�x�9���U�j�K�)�lTТ��[9�5'l%�ʬ`P��\��nZ�6\�0\	HO|'�pVz\D2=Xjw�$����TλK���!0c�z�0���0�$y%p�k