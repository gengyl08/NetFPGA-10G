XlxV64EB    4715    1250��7Pޘ�?��寰c"aw�^Ǥ=��v
Q[Y�̺"hʍj�Ac�����D�U���\�o҉g�8&N�|?�Q���o��>Xl��W4
Ư]<�vu̍��4���%1�T�MZ�O�<O��v�i�c;�F;E�̗��@U����nJ(e���C������
���9���d�j�j)��eZ��Ci�����AvD���-!����	������n9E�X��Ƕ�
]z��_�/h�����;�u74U�{����ϑ/�����
6g�[m*�g�g_! �����@ޱUw:YJ����9��[7�����/��-���R=WxY���e��H�c����ϋ�F.&A�(4�vd�7��>��g�����?��1� �DcK�����z�V�v�
�fn�D�I��"IJ��'Ϣ����}g�,�1�Af����7&��`��䤋��+=�(��^o������g+�oEk ��$��],9C)��e�O4�6�}Q����� ���ؤ7s��>�V2��5y��݁|�S�b��ޑ����1�1����AD���� "����O�Gg��=�6��T����NS�)�R�{?����cti��pֹ�����Y
[���G�&�F��C4��`�N�a���oxc��$��%C���d���S]�p�h�^H�P��_�S����y�EN��\�i),]@<��₩cê����"�6C�^��ğJ�u-���XLw��\`�p���5��5w�l�'�_<eL��3�yԏ��f��K޺�F�j�;����#�[�T�wk3c�Y�)��O�Xrg%,ɇ
h�����]1���$܍:&��R��¿�f<r�o�HE���E;�� �ւa��h�s����貢u�,���p*8��(�2�d�-hQl���4дIW��*C����&X�s}��/֎�?��@��Z+��ʡ�K	F��~�:����.c
�;Y;[�F,������[� @Z����T;:ȖUm���_�T�qeʹ���<nҚ�2cp�4���VC�I%�45���7��
Ϝ&!�N1����%�ç�5m��Y�*4��{���[ɡh�.�$��/���n�B��e|s��t����ـ�d������yI��)!52�,�Y�M��UEo8*�}JBk��5R ���= �,���R�|��	@�)��48�����>�H��&��Oѿ���Ρ��@��ƅ�}���n��S]j?�c	r�y(z�]�p��X]�(��|qV���.�����Ñ<��cB�l�awz��Ɣ���A3���gh���	�E=�V�e����&Ph��tl:x[��i5��X���g��1��W�7�_'��%�i���Ԁʽbz��*m��9WP���	";i2�D�7-w�T��Y���L$!�L�L��8aA�����y��E"j�YY�{�����F��H���}�q�;����ܖ����r����o�K�>t�&<����ct�ӑUI� jF�p��Ӱmz�R�3�t\��r��ib����X��-��"��W��w��tg�pʇ�y�^0�W�JK��z��/����D���p��o�-���I�,>W@ �񅋰G+R�k!#�CR� ���Ee�u��+�	�$���ȇ}���ЎH�����_:�=�|-�hJi��<�DxR��]��ֲ�2`���	�iK��	]�9h�� ��5jzq���� v��UD,J3CF�W�{����I �<�R��3P\G��{X��)�R��;����^�9!�6��"u�>]Q��5�Um��b0�gGн���c����:��A������T}EA����K��%��8x�X<m�C���b�W[xV;��`@��ԉBvMp^,��-�K��7���s����^�i�;v�C8�4������=?������ !�;��E�p�T��з����E���Ӆ��}kB����U!�x7�ېVI٦y`�8�I���
S�9��
]��T���g�yHy"\	�#$!	��I��C�u�D���PKV�#0b0H
O�I*�ѯ�;0���97��Ŧd�a_�y�;�9<�KD"q�����G�*"X8������ҋ@?b<����4�r���L��N�/Or�cc!,�U[X�P�'�UK��м<7rF�N#�::ώ�r���Rn��}�$�*�JM��Kn0~��\�f��{u����r�b�5����Β���2c��Gl���;�Z�	J�+�a����>��q)
ⴄl4�k�q+��
-/̓E�%�D����i���'�K�`��e���mzF���(m�RVF�a�`V
�y]�o���65_�u�M���O9����:���`F ��Ǟ��qYap޽���5��� dWu��jK�<��p�X(<�5{+=o�	h�"h
���h�j���*	�M*���oY�'-
�;�$r�ϫ~Sex�3��"¥6�Q��J��Fz�P$Ѓ�п�W0DC"�Mɩo��'T�Y�S�^�ۚY���	dݾ��ÃUo7���t�}�޸��ŷc|k(�amϝg����3NaI>�׷�UN��h���-�nh'(w|r��?gFIgE|��t:Ij4^*��v�k��XE���n-G����5�`���[�|��K�S��O�0��mYK�z���GE�YF�|>�o����b�?�m�5�@�t]M"��u\N_�@�v���oIm;��5{9LC6yU^iEC��}�����mc�Ơ*H��A��^��\I�����>Z"��+��n��\�zڑ�n���A�πR��9�/�wݐ��qD������i}7�-~[��>�"]�7�C�B(��W��n�5:ϫ�2řBz���ɂ!�춂myX[��֭� 	ܸ�B�Ż&iN�|���
ĝE�&$b5��g�Xv3Lt�Xtu:D��P�eb<?{,E�1��$ �%�ao��|�1�t��
�:�y4��F���F�=��3����i�Z����-��'��-��K�<��˭�#d���9x[=\g��&=���,��6�c.��I����	'�<ݬ������m��/��zJ��:�~+�t��~빼SrL�<��.g�Q��$�5���V ���A�^�A2N���e�b�c'AL� XIj�G��wqb�|[S�GED9�#�R���$��me���~�!"~X	mlz����Pf�5i6y۾A���BK�f����qfL�B�ְ`h��hf���/TY/ÆX�e��@f�K�l�+�Y6�Z�`Kdt�M;���=���XS���_��\+S��ee��w%��E�|�-�@Quϙ�%��9� �@R�ʃ��Ui�����oVL����~J�Z�7�H��IJ$i��M��U��A�����@_���B���"A=Yx׽v%1�����{˽5}\�]����hT����\o�Q�>��T�R�px�o5U�'~e��9����V��Z�Bb:4��R�+�3�`t��>	���޻g�F*������ p�Z�z����8l"�%\���W��[L�qb���O.X�����g�G[�ùz�;�,I��5�q�ѱaoh���}�+�k�>&�Xt�Χ�V�-�/�r����D��D��y�g:��dS��k/��,<�l�ֺ��s
SЦ��{"8=?נ��paA)�Zt�}J�����( �ط� �~��S��L���o_�n�{����P��ϵM;Xf��c�}$O�#�L���t݊(�ЪU�V9=<MN���+���E����F����׎���`���L��V���O�Z;.�Vgjfkr=��!���w�&���xtH�8.LI���d5$�@)�4d��(~��
pc�2��3��\�T$�	M��e�@��t@�P�j;��x*�i�{)��?>���X��A���ix�1$���+�d��4�a��t��=a�D��'q��Y܏���� �:�%��D6F~\ Kێ�!yc����ڔ�J_�
�; tZ(��C헹�z�<����mlओ��HYY�R��)k2�難zt_莽?���R
` ,�|ɺ��#��~����䁵Ϻli���Ӓ0�m��튒]��eQ]�q�E����fLb��G���΢]O�Y��w��y�x<��������˚�Z��ڤ����Q�q��3K��$Ť���Ba�����J��}djA<�K}���+@���CIج_�2pXQ;��_���A�&�t�1b�r�����o��bϞqӀ��4�!-+u#\�9�Gmu�!�eX���!yEAm�ts���89jZR���,�5�����43�Y�gP$�v�Z�'3����=�DX�lR��������3�'�E�Ur������}�a���oe�'Y������.>���SK"C���_���C.3����p��)`��G��՜nY��L^�]�_��j)��B��J��,����ٻ��`����ﬁd�����O�;����o)�" Ob��0��'R�f
8j�G�ܬp�t����]/�z  ��vE�?N��u�fx��WR��v��g-�5ԫ~�����,7�8MlM�M����3����("$0��h�"�A�!��R",!�