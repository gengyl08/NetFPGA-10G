XlxV64EB    221a     ae04��_�:�Kap��gH2��CL@n/�P���ӯ+T�욣���Y����x�R��K�-�-.ǆ���?	�Oc�w���Nf<�N.>�5Xn�l��^iK�y󢂀�Z���p�� ���(���c�+j%e�jl�X��m�u&~S�p�{U��Z[�l+N�.6�Ɍk�F��h��^8��`�Ŧǐ�5K�u��	��k�Z|��a�@�L��XcL��ЙL]�/�BY*�>=�O�7Z�9�4[s������l�2^����Ӧ�K:�uJ�ٳi�����+A_4iܓ��i�	�:V'�m��t �"R��n.���T���S��b˱Q��F0�Sa�������K.2�W�J�l����1E:�䰢z�[a�M���=���od�u:�u�(�T�ͷ�խ�L� �c�l�ҧ�����3Z��U����PuO�=6[�2���m�e�j[Η})��gz89g������Y�DV�Ҥ?�A�cTo�OoX�S�������\�9^(xV-�4���sB�-7�P!�qCS�1A�"�����֨��|��w�]�m��7BϤ���t������O�>�I��aoax#Q�}�w��~���@A���� �E�P��_���<��������@�'C���R2�`����}�\��5t�i��/mu{�G����6A(Қ���O/^:H���p��q@ӷU/�l�,αX/Ē�KM�uL��@ИO'�{����n����a]k�����^VKD����@�'�>��J)�^ �h����3
�$.��|H,�=��G �t s�@�"~�X��0v�܇/h88��a����s��j[����I�G�7�p냫�:JB*��͛��j�����r��/��3��� 0ǫ�� �=���æR����CC�N�7�3$K��m�[�O���`�ΝW�hX������;��D
�:��%Î>�k��E����w�ĊB��Rѯ�)���s |T�|��[5�/ҥ��G)��<��`����4�%�4q�ۇ~0��tտ� �n��-G�ң��5�)��n�Z̦*��ŻU��:-�~���m��%�	۬W�Ai�2	��<�֧�랮m�����x�3x\�����%�����Y��c{�A9G����z�O&���Ȭj�@�ܡ�&_����m�0������ �u����H���O��+#�I�~���ŕ�?��	��o@�1�mh���DZ��O���U�ڝ�L�j�_�\"��Ҽ:�D:�S=}b9�jP	Y�@3�C���4b>�*����S-��������r��d���O�X��M|��]�f��2z�q��*����.�^H�[��)����Ѳ�Z�j!B2̏�3�|�f�i������ľ���
i���TNp�Ǒ'���w鏥�~#�����C�A������]l�<:��s���\2��T}�:��C�=멮�ڥHj�C�	VH�@��Η����fS0����7D��'�@��V�}��U'ؽ�����+#ݷ�|%��1��T7I:t������{V�8?�3��)�o�:(J�&Ĵg��k�3E�&�`[�0Sh*)$��/����)���yJhq������yS��W��ԌN���z�%�$���Ĕ�ǚԗ�>U��MNO�74#� v=遄xSuʌZ�U���~�:��K���q�}���y���"���alU��R4�����y�Iʹ�j�8��`w��uH�/U�55�8bp\8q�:��s�>��B ����
�s�iq�a��:��^�s)Y������r_�X#h���pe�(
}��ڣ�9���Fđ�p=� DT�:Gy1��2O��ؓ�d�8��* �����5o�Y� F��K^�K�t�-*1:�zz��F��s�?�!�Am��G@�Q�4��0��Mh{���M���HMӑ�.�O�!f´�׵�lΩz7JY'Ϊ�KE�8\���U�\=�ٮݵ�k�N�1�9��3IКg�^�=�板.��r�莉�xB	8��7}O�R�k	2��c#F q��0����/"�꯴t��̸NG�lӃ�'(���!��=}���@FS-���UHx��:n@����&�{EX��j��u`UC�����C��Ǐ];�C�+���*)c���M�XXE���?�$ib"�4��d��l��\�L��5��=�a�C��*/�O���|�cW�U�4��T��P=u}�ɡ6�.|�[@v�ϪA����@�=�!���y[�U����˦�(�(v�/Ͷ�#�Vx�	�:��L�&n`��\�o���	�e�
��:(kG!�$r�_a	�~����o�b_11��[ɭ~oi��.�P~���}�a�2=��c����"�Y�y�@LE���G� �@�/��M�0n�A��G�<l�/�rI]���/YE�d�#��,�������-�bT��YO�J����u�>w�n�MF�29��_H|-$�+��U�C�On.`����\������*>�jz2\�tr�;HY�-���g��c}F?'k�����c�׆@�.�?FP������$�D&��V�Y��J_cY����`��8�sK�.�s�)혬]c'B��=ZG䣞+�τ��{3N�Y���ˇ��1֜�>l_�MQ!D8�:Y�h�i�n������$ǳ&<���-��V�g�: ��h?�,k�N�4�ЫTտˈ�^���`��J߬��h��Xo�l��h�8�)(�O.f��rS֚�b�(����