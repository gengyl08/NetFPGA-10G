XlxV64EB    fa00    2b303�}�ӯn��=��w����'K��˅�~����d��u,l�߫eD8�����\�6��g�EQa�V�{��Ո�盦Mwƨwe����(ca����FL��JPA��B�#]l�.K�yH�
Z1�Sw=--^�9*o���^�w�8�s
P�O~��IK�@m����y"�nDu*�'\��kZ:�n}N��ƛ�Q��Wޟ-�r+�V��B��N�9ѯ��� �Q˞H�gq'm)1+�eL���}U5c/�-�ң�����Y��5��b��?�yx�O\ �����v��X0���2LnY�7��W\����y�ݶ8<��p����>�/V�l����P�
vjQ�r)�z��6��Do��J�����]��Yg�x���r�)y�W]���`�����8�H�v-���,l���"a�h��*���/!�%U?Ui�>f)�(�N��x����Y��Ќ���ED�87�1��7C�(e����Ɏ6[1U;���`�C�N�!�9Xqm黻v��S׊��+!h�"`k�U.��غ��øo�{�'R������3��7p�_h��:Sb�n�F�?�F�����p�|b�)�;��d}%� �1�����6sD~�6��i��/gD��Q�f�35bɀn|�(,�G7�3| �C{����\ژ/|����{�!�s��Zt�M�[��@�}���.	I�B!]��
�z��?���&�:�;��/�1Q:����q����E܌P�1��\T�	/�11�J�2j=���.������F"��^�:�`�4�B����HzlU�uegtu�w/�}U㫸�_�D�|��!3%� '��iR��H��IЦi�B�ÑmA\�m���HѩL���L̡�d�Ғ�@"�����y��Pe)��iZ��\�K�闝3F�`<�2�P�2%(��e�}��Ԍ���q״�;`1�T��"^�3��.���ߕs��i;�l�k�uouK�/�_�/h�!��= :QT_^���)(:�Uq@����=��Sq���i
�hW�!��Z轢qW��	A�5L�kc(y�y�{.�`���`s%���0y�xs��Z�;1}�2�B����5BA)�/?~*��r3z�_��?�R�YM̭8���*H�?8�����G��O��#��p���s���f�P�S�'�W��"ʴ@*����߻lu��*~{h���zu:ᴶ���$��2���{�Z�Z�@]2�wJK ���p��|�wM��1GQ 5 �1R�+o����YeL������3a�y��W��l���ZN������4�{��$l�p��b��Q7{��"y�a�"yhJ,�9�V��P%ƀ�1T�]���a�LyP1l�7"����<�;
����WV��1��?4��_r��.��.�Ϋ�ٟE}2_�F�lw�M�6�:��TJiko�
�$��:;��
Ho����cj$��{p��z�gY؋�����k(Yu����hf�qv�0���(����"�Y~(����Ì]�l��t�o�9=٤��M=,��Kv���'���?�S�.�<�����p�]<`nƔPj��~�G�P�G�!s}gS�m��F�!!��`O� uD;�u�J��{�����6�`y�PW�|�=8�Ңl�L��\Uq"��0
���Qw`'���:�^�CP4ܓckM�(2���'Q(F���NUK
��aN����<Y��}���[:��E8S��x(��D��#"u:�@�_f�^��������&`6�B3+�CT��9W�Ȍ�mD֗��r����!,�Y�;����8�Q���x0a�/��[I��7+K�{|�u������D��G=Ɨ��I���H^nϬ
<N�
� )_��y��O���0s��$���H�ў>��¼Z���x�t7b<����T/�Jg��:X��w�^�Cm�諮���ݝhԾX�_��Q+�xߨ°����$���;�'��@��m"Ǫj�F�T�8~�U��j�,
�\��Ց��c�|�gd�(�kX�N�_����deo<��[k�F�tu�p�x��|?,���B����� V��1_�l��@K�{wQ��	�=�����[@��k
a�W2{��d\u��v�Y�ƛ�w(�����sN��l7�Kə�U3�^�k�\ԕ9����ڟ�L|�BK!��h���h�ڍn��x���ɪP&�MR 3���[��Or�]�F�N��}�Z2k���ȧ�� s��9lJ�;j�T��-&~j0���ɤ�m���g�뤓�̜갛"G�=T�a�?Ó�H� n\��F��V�Jfٍ&~tB �W��t\����e��P+U� eIQ��S4�;�Er�G�ko��J�UG�?+@d�)�FL_���<���vm)�E�8��3�p[�d%Q:�.	&i����Ge�cv xz�W���{�wy�%/����y��[:ݍ7��d+/��B?��k(�_^����;rYۤ�Z����Y�8�on'9t��,崒S������&�l�����}�eK���h���@��
$�$]`w�o��Ow��]�ͨ���Ɵ_8�nY�h�s�jnI�-���ru�%YY�����M�-��^>,
߷fvw�1։E������M{k��%�������x?}S�U�0���ft�㌾S���@������Q�^==�91GI0a댉D��t�Ȍme�g��M\��:v�Q��G����i/�����Y����F�kJ��dF�$B11������f"4?cƟ4�P	����Z��"̝��rK�fóx�c s�3.��,��:A����ij��,T��c�ɟXc�:�۞�F�u��tc>���ȗ�����P-��7�n}է��(���:.c���?���"���*pr�dWWӋBX�h�^�3�BF��r�P<���q,�;��̐ā�kKG@2턘)�|���ޡ�y!1^ҏ��t^��r���e�1�nA�D���9�w5�p���ݪ��k��J��zO�_,�>9&�XX9�s��D\��4[�*"'�SH��E}�����J�dΰ�[���� e���n�cIA�AՈ�?��6c�3��u��V}sn��+k�&Қ��g�M��-<��B!�M
����bO@����gL��y��Z��\�;�����N��H��֮��P$j�v��jm��ė��[��n<�s���S�vr(Q]v���;ߋ�N�Z�>̋z��������:�$��*2c�m�}1����^��~�	�x	���>0U�W��g�� ���+DW�q'�ؾ濖!*�3z�|�^9��x�$3.NV�� �k� �_�]��3��Ϳ��.z�ŏ�4�rE�qO����z���ǡ+k����ݟ8%������k�WB�
�^����Q.H	)��T�(����Ъ.ɖL� ?C�
��kFw3��)^�FȮ;Rbg�x���qc��GE���9k�4�!-����n���R�9[�'M_�$�����=�dV�U�������\���Ke��'1�z�B��'���E#���ڞ��u��I>�8��_�^��
��f�Q�pU��o����R�P�W������j��2T����*�X��o���bي�~IO����Hu���Y�h�ִ:�H��Cgq�K_�
r�Q�}MYP�3w��]F_�V;k0;�O�3�@XA��@�А�o�Y��Ƞ�ɩ�A�/aYS�,2ĸ���O�F{ƬшS�Mq<tJe�`6�=��I8]�c�^;�,Xu�0��#]�W'8{rt�Ga'��Ss�u_}�V�CT���I]kRų0B�D�ܵ3�e3�\���V3*utE�Vt�9G[?�6^�r58P�.|�]�IU8.�ɺQ�h�
���/+^t}*f!�@���'ˢ}eH/�g��z�Wj��϶�n��P���������� W�q+� ��:�I)&�4�Ѕ�(j�Ś:�����Pe����3i��ûD�5�rL�V
�4��A�F�0D�*�ppV��*$S�ۅ�+��H�qU�������X1��P7��=Jz��$4~Z�[#�V$�l:�W�V0=�@ʽR1�̚F���)�2~�q����������l0� :̯Ӿ��:J�(�v?=�*�����YO0�AR��u7���N�sh�NeU�^^t�@Hu��5j��cQ�i_��}��w��ƹ]���.���+���֯띛J&`�>�`Scb�$]x
B$Ih����JV{&��v�z�"� ���e�n*�	����CÄPZ��=S$k�'Ho��o"
�<[���=�e�%c��]�Q��*�n�K�-���n����󭴐E�ig�B	��n)�L�AL��N��֣5V�$S�N�S���\�c�R��7՟��h|W!�7�l�,�R2 -�*v0��{��eՈjG��:�~sz!��������ab�p"��1��]�j���;�KU����`Svq�\v)�lj\�,�V{wjő��&��ft�#8}�S�jz�=)|Kj��t�����~���������������U�E8}�d���tl���)���v�F���+�n���'g|��C7b�E�«,D�d�ī>,�,X�I��Ѥ|�&!/��Yjʅ�ހ�S�$���֋����{^�^��l�}Ա7+"C}j�ɬ12H��ߓ��U�U�R�^"���A^�_�aAҭ>�D��O���
W�p���������m���9�iG���QԖ�b��ŋL��n7�_����d��Җ���O��+���c��Vc�����P7V�'�	g"-�r���j4�EV�5�
�>W9��8R���iA^�) ���DB�G�ro��<U�i��6њ������EU&(��!-�}��zO�c�:]O���9�r���\�/P���B\%��mHpu2�5&���t����(9���zz�G�(���Z	�$�^+U��������o�[�
��n�#*�ﴗ����fF63�S*���*V�à�.�!��((J�f̀�������漹�AF7jD�Q��@zX$�r&#��g��쐋ր�F��P��q�c�PF��u��FZ8kB"����g���ly�7�� ;0����>F�w�h1P�|�o�X�'��H5�t°��5�6:�������)4��N��( ����YABm���_*6Ξ�5�|�޵p���(�4	�r�ۓ�k�l��}�bh��Pg��NZ��|.�������J�^�]�H>�QY$厍`X�~ӻ��� ��СVE�b���	/`q2�\�T.�ٵ�\¶��-X1f�rgM�!���w���"d�a7Zi���i���V�F�>	�w���nɏ��!������ER���8�p�ģhfn��i!�g�����?h�nE���ʇľ�v��^r��o��\�܃�3��}��u�ڶ	X�N�qh�
��*a�8L^�u�.Q��"�lf�9L�l&��`���qUC�J�TI�K��Eg@XZ�5I{.ƒ���,�(�Y9�!��$>9�t@ifk���(t'/���ںbL�	��x��(�B�0}\B�m�]�Y����p�D�A-�.�����ʐ��d�(Ȥ��:/��2c\δm��+K1j7�D%�^��4�P�{L�� ��6f�Ph?�<��T��@��%<U�܈`��,��G��ߓ+mN�꼢�2��Mk18�7�8��1�F�wLx99��g����c���{����yWnf�c{c<&#�+5bZ��j%�͌��IN��X�S2��c�u]_>��[��c����ܤr��\����:E����br�V�?�b�e��Ç�\�c�B5�s<5��X�T�/�8���<���U�aR�����~w]��]}�b�a�������
�8+Go�&��2������//���@ڀ��x�h�b�3��e�d�n@W����g{�8_���W�VJ���Dp�dsc'��4���
Jj_)� 41#I6������J� ��hB��+�^���ba:�(-Γ�KIA��H�"�B��H�H���!�A_�&�0߅��M�����d�%\�n0W��BB/������G2	r'#���i A;��=Ƹ*��q+�^�X4���&�\3��5"��PLu��	���D�K�<��e![�U���`)��Hx��dm-��;i�-���*��j��g�mf�$Ve�.��wW��/�K��e�W*F�y#q�6�-�}��֗G��t�2�;���u��hcY�̿��\��k>_�F�vV���4*���WM���=�� �^�/0l�na�d~���}��c��V	�C�ev} et�x�.x�r���"�=�W.9�>��ש4Y!94	������L��@~<�`#�9Z��)�f�<MU,n_�aiG��m<X��(	��8�Ԫ��~�Q�'�g�����9ϴ!r2���ɨtm���$�u�t�\�l19��E^�5��k�IWD'��x���[ý�{�E>��CD����o���m�Dq)H]����9�y:��K�ap�)Yi�)��V�.��'��4��ą��f���Kǉ9!Dgd��O*������Mo����H1�SǱ�
e�UxAZ�o���&r�D��!W������~�z5���7gl�
�@7�8��'*!�B?@��~�d��E����_��pK\Ţ��x�bkfJ���K��,1��rz�
��ԋ{�k���i�;i��P���ⱘ���OZC2��k�.�e��/I-T3,�zXݳq�M?���ڱe}�*Ľ�y\J��KI��X���X
�9��nd������I�7P����s���U����L�^d��@L�$[�)ۛZ�ӣm�Iv���w.f���j\�d�P�1�`�7�[������o�k���j��T��������b�XYDQH�<w�1ʖj��u�H1�<�@��h�?Y�S��۔�6d��6it��l*f��X�X�V���D{_�K��*�2.=���[�+�s�JƊ�0�`�B}��i���"��J=j7�Q�
d!��ط�/T9-����}�)�ŦDۇ�;'/��P�ڀ�Atu�h�L�݌��8�g:�E~��p���a��D:���&Ϫ�)2 �TTVɤ @�>��{}�͙�֜@uQ+�o�B���nNq9���@���#ֳQz9{,OX�}^�X�)���3<:��A�e���g�fZ���)��+4@Ҽ.h�e�0��;�
v]�]�}o�3��(���cwSL/��d)j^�+g�[v2s�)ޠV�K�D�H�ʜ�s���m���M�y 9���Y
�m��A�$���Uf՛��^T��XX�9�~�#�[	@�J���}���J]�N/��l��%b��aa�q!qU�i>^g��*jV~٥(�c�Y A̙:�	�)���ޙ�	��j�C,����;N_]Q��!�R�oP�l}c(�*����_,C�{?l�0�;l��)�Ķ�W�{�gw��\.gcf%k'����&�2�X���������s2�酢��ǈ�Q��09�p��7Q��/$�)J�[��:/6v����Q!L����t��1�u���_%S*a���H��Z�.���e�U��[���	���|����%],���D]L�h�%8C_!]�tg���k�Pݽڋm�[v�A�G $�Փ |��׾]p��d�`|Z��+�uܫp��u�ܪ�����UAF�)�E"�3�	vT'n�j�$ӂo�N�C��{�X!S׷�>��>�Pa�U ��Y��Leq�N�,#I}���h��S�?(����́�"ɀ�?>���J��)9�V�a=�꤫�O��A����Q���a	�c.EWD�\^���'�3m<���+�rh�U7�B/k��m�jD�؂��b��YZY�oz���tƊOnG^�Zfh1�8�J���:+����l�:Z�w+�E�>+Ӡ8��R�D��}���ۙ�Q�'�x�}��Q��f�Mt����ArP��~t/3����EG��_ɟ�1����};�!�r��Uq���ѱsY�������x�:�u䒯�"�EI�b�����ё۳_�QB�w���얱�>R�v�)�,�~`U�ly[ǠI�0u���嬕���+�v?c7\��8ܤ54!�#HPma,˟�fb7zD��ϊ���Y1���\u������W���2a�2����V��[*��g�<$���^"u/��������G�f���<�#�K�+o0q��J�c���N��w#�Ѷ��ĺ��{2����r�" p	����(��վ�����@n��_��b����� 4$�i�_4�ƌm��#��&��,��\��\����M�S�cfTe����*���UW�~��������t͇rvKh�}wX<q�7E�Wp�`�C&���D���M���D����<��x��S��Ǫ�T��q\��j���6OȺ������|$�9ᒌvdm������nH>;���l��� ��x�p��C
��Y�לLڀ���.n�%��&������]x�:�G��4_DRD�w��0�g��FV!�3"��~F>�(?)U%���2�R2GW�.=N�.��z׉<�0	�b5t�&luV��Æ�������'v+;����uO���x��2f8`5����Lh��\� :����L�<�\�^p�\�7;9&0 �93�`+��h���#���x8���r_7ĭ��V�6 0ݷ�9���Z ��5��gk�ΣP�'��5	�w@���� $����UM�ؗH�����fS&��xJ���0�b���q:&z|Ej(��cU�ܐ0曣bIĘ�.����z&;�l����t��0$��(S��xY��������#L�(u/�1�d������b�ͻ^�k�<��I%ys���L�Q΄�0xL�"��޻d[D�!��C���ά�?�[$�k;�eN��jz\��Az���$��!�N�6RX%|�ⷧR�F�>H=��Q�7ԫF�͎��7*S$��5*��
����p枬R<��-�@,�
��(�B/}����m�����8�ɒt��	1e�W�Q���O���)�o�6�_�sѮX��s4Q����s*g5����G_�ǜLI)���:�%��^*E[�����Z�x߂�|�Ν�w	����E�0���LH{Ɍ+�O���\�P+��zQ��BP>�"c����q-����TA����=���<lt��������7���?�4T��:Zi&Y}�:���eK��|.�X���$�������m{
u��̈��/n���Β9�94�i�S���t?%�_�d�fɄ�P�̩f�ԁB��S����i�y{T3�;��e���Sμ@�)`��ܗ/���־�!�?�j�4� �bi�{5f��_I����L���ko.T�gA/��͝c� kM\�$�\���.L���-��r.C�H���~�x�V�3@9��E��ByC��(E�_�K�5�%Fx⎑�L�F���ݢ|#n���R(o�ҡ3*d6�;0��mB&ȸ�&~ʄO z������Z'I�i�}�g\�� O�d_qq6���1��E��;���X��wA����)x�w�`ｫp/����J-ܽ��q>��U�p!t���r����f���o��MߊY/r��'y*
�#+G Y��0)��F���P���8��y�&p�kv�p�C���((�tN&�fG���L��NV�)�����»�Y�3��{��Ė�,�UY��k�$�ZD�`�-��g*j��g�a>(bY�A����s(����c9�C��OB(|����;�Xȋ�Yc�H��ɒL�����v���Zjq���z��a`�2jO����he{E ȍJ�KC�n �~uTR��jɻ+9c���e���'�[\�+�S�#��!0Դ&852�3(W\������S/P����~��;�s�8��|�F�SOs�Z�u&$=&�R�w���:��>4��n2$9�4�q+�є-�v���G\T�Q�Bv��ti�TGT�p�e�@2.U�U�|e�a9m�(M�F����ʗ���v�~'���7x�Q��2��Zr��Y}����W�b�jǈ�{n���N���2TD������	Q�`i�5�nDz��}.�J̱��h��Gh��B@{�?R9%v9�ǯ��B-�s�s�[�c���W���{�b�׀�ŌTl5�UB���"��`���nɷ,BZb��Z�ua�	g��.���vA�����)+���q�����t-�[�����
�(���v�Y��&��<������=5�oH|�[�\�W;�3�-��n�a4�T�Z�M����EĜԋl�����!�x�z£�|Lvʁ Ly��?��d��*�h��ң�:HB[�ω��h �$q���_���R��b�C�t�f���.���0�~���^;���u|�wU�&kx��Y*���S�CDgD��q������I�a��۪��R+//i�y�wh��鼚;Okf=o�k���%�b*���9��K���?��k�yڧQ5`l��Q)fp���@3U�wzL��~��P��]���+�j���t?w��@���D���$����m�X���W>ҽkOV�~�3(!"�SK����\�'�
��$���7/�2�/��0�"�q~�M����B���P�Ƽ"��r�-1�z}��$���vO|����ir��7{+!��N�1�y�ue�z]����䲀�l�.:����#�ݺ��M�Z�K��q��`�s ޿�#C2\j���%S+������� Ibk�KILu$M�A��nYE�g��Vjݶ����JÖ�.� q�Zr�`&ه~�
OZ*4�<���H��j�6�i�X��r,�Q��]@�уQ�s�'J;�B��XlxV64EB    fa00    27c0��s��<��6�[/�ul����(�EV���Q�sơ"�0��͖f^6sG�ݐt��
X6��:�h��
�Q����P"��i����m���4�o�Rך�,��r5�޲�W��;�*,^CUnx�A��Xg�BZ��
 �A�b�7�0���6�7Z�g%����6��u�:�{:��+欨 R���Z�+�Kܽ��3� ��,�!�H��#v�S�	P�#��6N��~Ć�Z$�)Ra^�X�|St��l�T�p ��"�&y2�"�G�D��UGe�`����簲�< �:7jc<�J,�}�fk���8 ����+���G�LTq���7a��� �W�	�qN8��Ew�\f���r���a)�Y3�3���M��h�T�Wq
�
�:2����ݟ[~D�7�Z6 /> ͬ:�}�����m��4 �3���P�Wo4�tQ�t�%�S ,0!��c�;o�z�r��������d
��s�|#ܛ?��,|)qs�ɵ�a�J��#�������'Nx���_q&����2��0�{~UW��3F{x#�֫iE���RGÝk=�z��'���EA�Ç�Wu�W�>��l)��6�@�W	`#:F��Ĩ����e!����P|��ù�K���� ���ZN�YiHo:�:����T��R��mD�x�B&4Gc�[qOKv��S�z�`��l-����HӝqSH+d�#�s�m�NrW!�]'��c�eZ��D��4��P�dt�w���.֗7���A5k�K�r����0�u�o} h2���)ʅ�ѧ=)Vl�Nò�V�ShO�PY!�>Ʌ�[�"������W����7���t`�As,ۂ�n
w��.�����y�����ct3C��Ж�����>0JG�dp��Z����+P�/����0����ЧO�n�c�����qxk�^�l����|��w���s���\-�16ZC�P!���,n�yU`�fՠN����cf�vLVǪ��FqҌT��T��s༝^\;�1�ެ������Ҟ�0^�!fq!{dU=�u��F��r3�K��?��J��:�0��Tp����x�b��R�L���Bhd�0Re@yxI'g�ؙ����D�*0�q.��5>�ڭц>�ڣ�@P(V��~<Y"`V�q�&��4��1����B���P��xY���o�x�a�D�<�S�#���Y���(M�|�f$���4������s��F$�!/cE�H�
q3��#m����C��+OI+ !��o�}c�� 5�:
W�}����ߩ+��� D�~N�D�ࡋ?�I�fX(����|��$ؐlo�:A�A�a�x�/�������#�k�C%�iGeݗI�uU:=�n��X�+t�ԣr1���Z~�N��J�)H򭠧ƮMk?��yG��.;�W]�Ó�I�a1nJ/�ܜJv2z�Tac�X�����{ɵ�B��nq��eL�O�_ߓ���Yo,8[���lG��m���q��;�#����}�)D[I��/�ާ���*�����Ouxi����Ut���uY�I���o��
K ���cC�OB�t�iC�>M��6�Q�����ا���OC���4|�	!O=o$�Lc��?�:���<18�F��-z��W��F�NV�Q��h|i(׸jꎻ����v�q aH�"����9�wm`��� ���,xd�Ԫ�FCEV�[O��Xl,X�pU7�g��'e��r�.������vqu���"?w�)�I���7\�����r2�]
�Y/*��ho#�	G��JZE�n�5���o6�Ye�����3`�Pt��D�'K^��Z%i,���Ԯ�{w�Kx(9;R��	��kP����������I�j��VnH-4��w���V����A�qU�4LK�z�GE�������i8�zj����v�#n��ЖR%�7F(���y�-/��pC��M�/�L`!.	��L��{��!�A�l3����4�֭���hP��bʋ9���-��<�� +3^�M~�o[c+�jVs5�υ�_M$6��BN�8k��;@˨���q�Y�~!�uN*�ĺIj��������/�4�S�yq�G@��ނ�鳸d��_�*x,ys2D�� �ϢSb s3@�
:��IB<���uj������<�N].���fKf��g�?!?:�����xb�g���N[Y����HD�0l���	�0�P	X��Bn��7�ǸȒB���~�v���T�0~+����5�'0ͦ)��Փ?c�@#���~�����j�3n�z�­�I���S�ҕ���]O���u�	IȖc�ᴧ��� �{�{~��#+�Y�*7\�(��B�
k?��K#�x�9 t�9��F�J����+a��H��9x���t%4/�����q��O]����S&�;y�֓�O���M���W�jؘ9m:��F�(����Sq�	_����5�ut@�c�]Μ�ѧh�� s/Z�����+�r �!ۣiE6h;���"����sw�ѳ~i���}�,y�����r`���L������('���(3iQ�OP��F[|��I@w��dq[`��<!�T5��eT�G��l[�Y*�@���3��(]@q�~	~�dr��Ut�
>S�o���>�P��������2�$5�=?Z��nJ5C{F� ZU�T�%/C�#P��8�RH�6Hl�����dJ S>�p�35[G@S�+@}��n�~����&0(�K�"�r�+?����5�(�j���\�f�~�S�3N���'��;�WDxV��>��;�誝�K�*ʹ\�j���.����oy�.���0� ����&����b:�@�PP���z�^�u��zl��m�������o���
�~�ݢF�o���@�-�
U�!�Q���e����Z9��@h��;�NT�X���s��v�*z�kd��&�x��9co�JW�~�dm1���D1��D0��3j�>�=��rb$�`��&�>z&���1���a?�����[$kV�bX�ҷ)�_��v`�E��<+�(�L�Ҳ
~z
��Ş�!������p�7����+���KB
v���3j?�f�$7
�١&+�%|n�{pI(�|{mU�ˉ4��B�$��#Kښ��?	�o��T�$+qr��ך/��>�9�nt�����7U��VD4\FT���3c��wr1����r�5bM6?���pN�[T�}�d7��d4���)Jw���R"�%����pE�� ��U� 9�qah ��
�����"|����I,%���e<������PS��;�e���%!�.�_B��+uW����%QRR��|��&��ޞc��֝RW��ّ�9��R�PZ��MM۩$-z���V��X�Ӿ�t֗��P?���U��!!D�}j�X͛ e�dG/�C�Z`��N܋�B=&���%��3�T/����}���]x��΢�
5J����S���D��p|Q$+�)i���8��µ�?�$&�u8��u�$��*�w泎( nT���A�ý��\���7}.�=F�Ǯq��4ēYߧk0>[.�]$�q/|1��}�<xa���R�~`8�a�!�g�7��u�˻kaR#�
�)����
c����<�Z��%n$'��z]�]���g��b)�x�x�E�9Ҁ�N����*�����J�k�}���&�����Cl�!�@MB%�	9K��_�A(�?�ɞ*|��L��%ld�+����σc	Y/<��!�חO`M��E�Ie�ޕ�瓯rܫ_�>x�M��{'�S�#q���lUs@�*�D�?�\W�v]h��8F}�C�<�n3����ş��<ҷ$nH>�U����y�EB7>̪ơf�q'|w�X;̱h�"qc5N�E�D#�V��â�Eʁ4�#e��QJ�q{��oX�M��\�2X�
��*�o�i�a�i
��2�p�M6	:��E��<0�9�,O�~�r��4���Q� $�����D�n���d+K�=g+8���bj�c�[�x���j�I�ⴟ�2	A�ݟbm.A��?�4')��U��'�6��s��#'#)�GZ�����֋;���l�Oߎ�c[K����)^�rP՝D$h��S#z�d0��)�j���"�r�����5gOu�z#�qֲ�ݙ�vR�| b3V���%ݲ���zK^8պ@18.uoɷ¨t~sZ o��?��b����>�ㅉ��&��Yk�Z�]�'Y
�酳ٗÆ
��a�-f�:;Z��c�x�^�f��P0d�$��u5�f�Q:�/�K��A���3/J��Ox���n��۴r��go������ޞ�En��v��?f��g&�B�G� sq(拗ۣ1�b(b�q�&�l �ʈ�������fG�lf����kO��F��|D�٫�-!��z��b¼��o��������>���J95 ]V�O|���Gd��i����O���̢at��O8N=�`�	>�t6��_����X����Osv
��لTYD"C
��ڡ'l��I�?���$��+M��p|w{��s��TU��\C���IU�@�N�q��$"~m�^,G��D�p:HMv,6R�P���X��e�B�[T�ܘ �������9�r�iy�o��A�W�`���HqŔ]�n������&������*�g+�!�d���-޼��X�X�d�E㉶�o�;����xo���Qӑ�PU�Z]v��|�Jy�q��%-�ӢJ�,��J�MV�(�Sl ui��R����_� d���EǁO���ł/���ɣ`��x5.�P���t�:�:�;�pQǱDL���%����bv�äɾյT��6���
�"�-wt� AMD������<^g�=mV`�#X��v�vT��
^�Q��m�Y� *�ߠd�T����/$;$v(��S��e����&+)M�p���P�6(^pA�z����X��c��Wէ�(��a������B\!x�L��,����
���zb-(�ґ�o�-��:�L$��H~Tk4�[�b�@���TǯU���j�2��><o4���u��]l��ũɭfmJ�z�����*<��\^Ĕ2=��ꔛ�F������.�ւ���c�D<��p�LC�gή��fd�-�󹮐K�
Q�4k�t����/��
(�H�q [��P�����ʍ[��b8J���aL+9d�	\��82�-dp��AIt���}��{?��h�\�!Ƙ)y�qh����x�m� ��VHD�/~X�ke	�	.�&�"i�Y�[lx�{l��eeA.�Go��㿙�D�Νmn�U� �ry��:��/�s���_6(��h9�|�FuaX�"v��]�����S�%�SU
Q+FLы:�Ꟑ>�J�tp���Epr���ٍ2
-�/M���R�;�s�?;\1���e:�,��93R=}�ɤ����W���ɳ�4�Bf��Ґ��+��+9�C�tq��f���h���O\�,�]������j`9���T���p�
WΤ�����vi9��wtI��q��>� �Y(�)f��ΓԊ��fp����-Ff�k�P����{�8?
�`��KEy'���FAD��C�^j�F����)��A���wiҏ���7�4���X'̉����u��^NO&����;LF��:�_���k�=r�r#8��jA��J�V|���	��7���_X���]��ޒf�UͫO���Ο�eθ�Rڪ��y㆟{[��3/̅� ��j-%�9�|h������'��2'[՝&`=~{帖�yH�]�������} �R$؜j*�%��|�6'�I�/��n_���fˡ2M�-a;�S���-�'%�?�㐐�3��J���-�:���v�a5�� �y]D"*��2��I��4DC���{yG٘!�`�5�"�rcX�}��Bƪf�-0L60�GQ�Z��^UUyI
�2��'����K��znTC�ׇ��J�>�λ:���7��i�S6�ئ>y2[.$]�G ���~��]�����j��c{ȿ" w'�W�_i�V�ŉ�ԷD����hzL����N��ǂ�#���M?��1g(f�~d�h(�о?uc�%T���� 0{���'�p[0�Y-YRF!;u�|Z�7l���2)W"uq�b�c�+��y��i�dG��[�c����"m�[6JJ*����ݙ�����k��Y�`gg��sy9��z�: �K����6wa"+�QKj�������l	2��A[m��^�hդ��O���P_�ɼ�-{�V���d�R��#�������%��n���WY�~���h�~�[+Y��g��J���P'G�$\~e�����d�{F���ꙩ�`���*$�E�u�f����!�4ܧ���vvWK,P􋕋tf$2D߯���s�'~B�����BGJ�0��q�0O�;_���V���#�����ԧ����Q�ֶJA�dGf��������~�9)A���w�N.��Y��4��&B��FbPs��L�K=*a��?m���pz�0��+�C3���$�q�L��\�%�-�;���������9'���u��
��j6���J���K.?�&<;��3�����R81��A�-��!-����0����J G�xo��c�Lz`��E�R�8Rmf� ��u��=>�~��BrI7�����_���#����_�������)T���h�G4-AK�#�8�����f��ր��w!�)Wo������V��oo�����?�ha�}�z�SW*�Օ9��,?��Z�*��	+Y����А���_S��Rp����*Y�B��@�<��
MX�����t{�_Iٷ�i�{2a������0
��F+�E�y��K�Ԓy�O��w[O��Wmo&�2�ؿL��Ĺx	���EP�r2���\���Kq��* ���9�`�-�������7@��*�e�f����Tu����I���u��	Nn����i�����g�=H6���R{�yZ䷥�B\@��+p�vN�M��F����P�|��U���ZZ�o�m9h���.?��s0�Oc�)�u;��H���Ӧ��K�x�f`[^x,ߗƢ�Q����;\�e`0����V��k-���2� CD�&��aT��L��H��#�8�Y\��F]�5l��P�m|a6C����u�+�?��s�Qlo5a���ю$l(ʝF�6���Q8���XN�`%X �ް��T����?k��7���ע�^cb%��?!���=���f�4������s��o� ޓ��&vI�{t�q# �Z��)�s˂4.�(}��Y��K���V�r	Wf��C����z�LLn
8�*<�������\^�Jѱ�dn�{X��[Z���Y���������%kԙ9/�^_V��a2���<�NϾ�& ���zG���O�\�B��X�f`�ϸ�ߎ睂��&�\/�&��	W���e���y�Ey��%d��Ǖ���{JT*ͧZ�!�'(������J�\m�vA�GC�X�JDWAݯ�b_`5�!�L*�� ���R�J��v�D:\��mSY�4����N��P�FG�_�KP:ZO���:�q��������{I��� 6r���*�(8S3�;tv�0$p���H@� C� Vw�h�������Y&!���dW�ЌR>���V��x��]$�:�i�0��I�֥�%) u׆�d�9�ǐ���j\�YbՇH/�����[��4 ��� 
ؚ9������ms�#͂��=ՙ�� H�ᇗiz�V��]��f�R�	�u��e���|𩷇����i�j�h�?����+t�c�d6ί[���c���`4�i���*����x���f��f��a��%�ȟ����Zg�qu�먫��0����=#&�o�����Rbm�ӐwOk�o����{��AS���d��מ�A��|_fL�;4��;�N�q�um'�o�6,�u�큊�^I �a��,��#������I4mYH�m�(�й+n�>!L��p��'��[2{�1�Ӝy�{�j5�&w��W
�sН���$/ t6q�C�DP���lX@Q���3���;
��6��`?b����9*�j��]P�Gڭ�t3}�\3�Do'L�I���b�lzҀ�)��P;K1[����]�8a���>=S�nW��I��.q���Pً�.S{^C^%�X�;��:G��扭���a͑���Ya��?˥�[?��y9Z��t!�cr�C\#�n=9��}��+,��PR�S��^ʜf`�Agf6.e% ��82I��&��i���w-1��0o%��/�9�c0���Cuaj
�^iR�v�R\��neCCb��cR̹ �{���s��\t�<��9�U�j?n`5��[l�Kל=V]zx5�X&o�s}�[����k�P5/[W�xbb�n�c"o�X�󞤴�{��wv�����5^�P�W��.����k}�2^NS�dK`��º>ew�����D�h�2rΗ�+�����6gq�Ĝ���pg)�X���zl�/2���e�zm^�n[�.E�]UK�^0��ێ��W��T�Ɖ�kw�^�$k�Mň��Pɼ��Q�'σCI�i�Al��j`��?���{�
B&$>��UL��r�oM�dy#��kNP���Xꪦ����{	���Qm���yL���^�����x�
E;��U�1�7`�	`�c�iWq�X�d?��N�s���v|��-�>�&;z3��I�b�_.�$�&�o�`��m==�p�*~���W�UKЌl���@C�ѕ�v��E
��p�X)R�Q.��Gp<�8E��t�ϵ65�?ן�
^�#��u�Eӛ}}we�I�5�)�۵��i12AD��q�@�K�w=NNpk�	ݶ7Fͭ ��tW��D$+WO�gɨB=c�30��7AL�r�2�h_�����o�ϊ9談s�"�ǹ󈒒t�=�{P�U&��i�+a�ӌI����I����nӗp�v��]]�IŎ��=n��;T0�q�#�2�M|[}=���esgv1J��<�JAS���7.�U QF�\G\�T��/%��(Y_eLt�70P��B�1"\�4�Za\�Q��<	��B�xH�!nN� :!*�d�����Ձ矍�eX+0Bgs%�l�AR�)}�˨�f�7V�k�l�<<��;l=n۩bGV��ӂ�h����pt�'B�������E�%T~O13��Hݘ�4�c>R�ڳ;�))��P}Q��ٸ��6�v�#���g��mO�Eڅ�1�$���-��Or���
��2�r��M�WJ�^�@ʢ�M��E�̀����F@"X�����fc��[k�8��g��ނ� ��G59��cK��y=�ܬ4��*�'D������w }�!]��iĺ�#���*����q�k�|��+A5ؔ>b����#�^��"���ڈ����� ����ы�s�s�Gc��&��%�J��4��9�����Z~��zS�r��$J�F��B��L�j P�}8�J�-���V�;�#���Sz��~u������۪����^V��9|My8��cQ:�Z��������õl+�w:�g��h�*�*e�-��+��o�N��p�Pd�8q�4�f�%?a9��C��&������Yic�h�ӝ� dP-Z��Z����
�4w��r�S��_������B�}��[h$�3Bk)�� �ހ����^~�{64��d�{�����	�?�8�M�f��)E��#5��l����j���N�B�W�h�(
��MO�1qH}��̕)4ަmp69L䳮�O7z��]��8>�(�o�zt�̽���ua�λ��=A�A�f�Ӥ��̸A��q��(��R�*�>xH�l�e���H�'�8�}�gC���):�o�Iq���g19�%O��S�<��'���`|�zA�m,h�1t�ܣL��렯yk�GE7��"���XlxV64EB    147b     500�������=J���:��P�&);w�A�YQ*U�D�٘}4I�b�7��r��"�skj�`�\�o�.B��v+���X�2�B���iV�������ѫ�6e0aBN�jNTJAFD�3�;�N������XE?����ٰ#����\f��-9�Cخ_���Ć
����Wy䥋��C�j�^�P�t�o
�'����L�3'9�cf��'���7�\���j������L�F��T�&!GPĀ��<X����c�\�g�	�S|wx�HVc3:��Ju�N; AK�jP��wD́P͌�jߍ��>1	���${.l��7"����^��ϡE�&qtdǹ]io��}�6l!��Oiu�n�"l.����-&�Q�f�F��c��)B#�b)� 5�Gt�`�V���:!��̅�i^��̳���?W�[����>���ӥ�g|B�?��Ҋ�mUj6��IL����é"���yl� ���{��ƜM��`F+�7�dD1����8�>���D�U����f�F�>�d&�u��A�L�����3�S,	��+��S�ӱ�y<>p�FS��o��v8���t���1���_F�˯ȗ;��"e�1ˉVS�cT��w�Q�vK��" ��Aں$�ݑS����%��ɴ�'/+lb@�U�q5���CH���0y������C�BG���Wԩ�u��E�ʪ&������U���kQQu�u���{�q�~-w$Ĥ�LDܱ{�������O2w��2�kԲ��Ǎ�� [\��j�`��UO�;�h��\��:�m�H�r#��8���#���ʌe����`���u5vIm�)t�E;@uo/t�QxP[��2oF5���޻�����F����(f�nc�JZ		��Fk\|ɇ�l�?��]�I����]7��ף�w����ľ��rc��!�VWa����q�v$ᾑ�M2�R�NX4�J�1�@��i�0����Mc�(J`6�~;Nr�!������I���ɒ���Vo�#ʺT�tsl�_�f-o�*���������`W&riB:0�M����:1��?�ՖW��';�ڛ��+`�p������rk��d���	ҦT�W�β ���9j�W�}�0�DT�W
X! �~F��8��N F�їW��TZ7?�������訊�&C��F%X��Ԫ�_��ݣT��G$
��Y��Og]c�&Ҕ�4����&�ӺiBB�U@�:|�!/����Q�B���[3�WM�