XlxV64EB    c9ce    1a40�o���c	���g�,5��� �h4U��Ple
i@�v.^��'�7+�m�� ����YQ`$.=~�$OP/�|�h��uޕ�r����cu��32�;�4����6䉺�H�w��2tk�*�	b1�y>��(�n+�9����xi�*�3�bsF���:����bl���)ɁOV���[�GQP�ZI ��E�]���4QP�ΰ�1V��mk���b�o����_Ǚ�0��՜F���r@	HN
�1��2��u��PI�#���- ����*��4(���hY]��t��9M��p��,���Bi�[�?v!��>6JrX���1y?[0&�������;�4?}s�5 �8�j��5��&�A�+�L
rD�jMkU�(��-5�J1�7������P��X�%Dy&*�Iy^��p�e$.*hn詞r�zv�Q�Ӓ� NR����|��^��c@.�}��J�5�F���Z]��)�Z�s �����S?&q��]d���9R���F�|i��r�hE���yh���ߗy�sb�׏��EB�
(l��z6'�NJm��X�� ̪���^�b�b�!��^9�1���z:Z���kiǘ�}�\,C�F�M~j�?)|�p�9l~`�hw%�� Я堞Hge��  .���D��Z�З8�̽\��\$�;��d{�E�����[�k}���T��o1�l��O��k�R1����BT�ӄ��x�N������ �E2��ºp���p`Uɦ�5�iT�ڔ=����Gc3+�2���D;v�U����"2�1�dM9@I{@��-��x��2����z�E�J�}6O�u�7�yw���F�Z^�Y�!V���G)a��I�w�aբ����<::L�)���D�m�r��x�]�<6�wT�ӯ�.>��CT��A� ��]p�
���9>E�^��c��޿�n�  �ε%n�ۃشT3/k0j�q_~�+/Y/C"T3��#l�<�O5���@-� dH��yY�jv�����[g��$-Z��{-����fk�#��)���9�m����]n�����u�]Ij�A�͆�[�l��B��Os�=�#:�qV�M�9�s�����Cᇶ�S �w��hS��H�C�4�����]#�-��]�wl4�����)�tbᴚ��ꑷ����.�ﱃ�ɒ�C���P��E������G'�=7���?6���t�H����X����2��9���EC�1�ޑ���KP�uV�ɓ0�ɶ�<|J��j`��37��F����Z�(@�$#�Z��=�cS�7��\F����_�}k,6��y�(���x`��M߇������I��|��P�+�Y_��$q�
�z�'�f)�'U)��Hd���%6
b�dk���mX����;gz��|���)�Σ�]��q�SH��u�6��ݴlf����G�ܟ�����*�����V��L�n���Rc�`a�����$�f"��6�A�D�$����g� ��7�-K�_�n*�<'<�Zb���Er�o�P��퓟�����֧+����D(��;	�t�B�\N�W����چ�+�W\������%T(p\�:���_bˣ���&`v�7�%����$���,M�^�=����`���`/���32�v�f]Ot>e�߃p��+r(qʇ�V@/S��դ��'߇��R�.��1��Dɗ�܌���22YN����6T�U���h�^6�/R����?7̀�]~�B5G�M�(as����2�7G�C�x�bԄ!~�6k��Q:a{�)v6�R8a�Z>A�W�6��ٯ�$��"-�pi�n&�`0&`U`��A�SE��B\��������9�f�������UQ\c�O���c>R��h�Q�9�-��WR��~j:�߆���k�9�q�r���r�[�����#P���Z �7>'�C���jz����.1D��f��^�l��0mo�/	��e��m�J��|ƿ+Ia<l�b$�ȿC�]#t� �Mm�p�GO�zFh��6���|����6�O���y��ʈ$��1�j;=�4g"�^�r&!��h�C��)���=��ai{�u��~I�p�݂v�1G�KV�����w@���}V���n������<�`�T�#�l��q;׾�vzw�dw÷�
�#DZh�E�u�����ЦN�W[��wN�͐l�*ueQ�&�Y:#��2�l���xX����w!(9���K��w���nל!2g)��U�q&;�/����އR�9s���"����
o��#��u�ƾC�7�C�v����V��.���Pq5PjPP�:F�TcɬZ7:{�*��5K s|����dȳ�E���ge�5e��/�P:�q�&�\�z�����R#�;E��9���b�?u�U���R�"�P�ߜ/�ĵ0���Q�ʇ�eU�{��ao�y�w@�К�$5��ڨ�A,g���=����{����C�g�i��G��l�@� ��뻣�<����W�acM���Za
��W�:�+�C�FMT=�Y��A�]8|j���\��]&׮�V�R��/�ޘ�w7��	��L��MP.c@l�&,j��Nt��cт�:m�Z�DB�_�����DZm��BŔ�7��ㅬ�}��E��〿H���}!�Cߔ?i�3Eg�}��[|�p�S�5F��\Ut�1�Ch��*t��e���W>f�GB�_? H���	$��SY�k%�cZt��֘��;�r��y�����!_ ��M'�b5��	l�+�y$���f���eU�6҂��X�ۦJT�a�&*�^�*�4H�����L9!X�����s6�5d�i���i�&�_�{o����q�X󿪱s��P{���Xߣ�>I*K���hC����͸�HcХi��Byn��{���'�.%�~��A �(r���bT����U�uK2���G�'�!�A6c��m'��SU_0�hD
��n=AG�N"O�:*��_8�������������Zk�C� ]R�z�^����O����>|��f�7=�'.�f��l����b� ���=}2�h��L^��&���S�y��N��r�%]�
`-�������\֔�����H,u�XU"�ا|�M��,H�]�-�2�8�]���wZE~�����)�Q(�^y�L&c"[+�� �{���z��Y.��욚��' ���f1c�N�%�n�Su�K-�
�Y'O?-QE�F�V�<���'Xi�PY��c�˒��JC�X_����#����MHd�*�wZy��>�r��͸�$h'���F��+�>�� O6@T���g���-�J"�HG"\�Z�ISC����ꗓ���01�4|��i��V��ަs���hFţ8�4!%#���"_ƅ%{�Y���,��>z�� @L�o�7���^�د���n�cU$�\�}��b�k�c{�Dl�!���d�m�������l���{0I��q.�M��R��$�&-�	�� ���;iŗ����� \���	Z�G�^�Jk�D�S�I�U!mj�W�`g�;��a{�+�6�	�1*_��J���=�_�H��|
n�L��O��c��"wb4�ݗ�iן�0���q/�����y:M4����2M�zá� �5�zx��ހ3J�w�
�h�j*:����%��<�Hk�!x^��A�����B�@�!|4�	#����棜 xqq�v������:��ΐ��&�-�Z�1=�ݙ�۝����hD"��5/�Z'yY�d��T�
}iЧt+��۪�Y;6��w�����R6o���Ӽ���
K�LW�W� ��h��קز7������7��)<\,b�z�l`&�X�dY-xҥ��d<
:��<�;M�#Sa������v�E��t��<>�z�Nb�B��v�M(�ֈ�M$��@��j��d����-ffuL�|@������ ��[i #��y:�,��WMD���Y�u띦e�nOg�I�x��yW��k�^�2�4�>��Z�ɬ���Ӆ�+��|3yO��0rf�C� ��Ș�CO	Ě��Ay�??]�H]�wՑc�y��}3@5N��j=���;�'e<b4��t�ʯA�ޞ�I�H����k��q� ii�TAz~J�c�}��^R�l�:�S�n�6C(h�k�^��k��Ta)�m�d,H�W9^�|5IF8iWo�rV^����'�v���gܹ�w�0 o�6V\����e(dE�V����~MUed�s؃Yv�D��gY�v�{/,�{�4�-O�&����3�Ɠ�ɉ�j2�6�$1��F�XC����x±�T�px�o>��d#�cՋ�	
��z:��#�,UK�x��=:�*�kmu�X��F���z&�	<���bF���fK�50dE!�5�s�e�%>x=����t��P�'XrvR��3���N������
�-TJ/�ZpӪ��=���&���}�)�'&7�t<�>�����.��������s�J���s;F�Ժ��h�@�ek���T�㞟(w�9,���$}JV	8m����tۿHwї�cש+�AЈV {�ϵ�t��w�����}��(�!�@�3��;��(c-v?��>���?G�_�η�6�po��D�FlBKyY���0t��BL������6j�M�%J ����E�82B.%�3"���gt����zA<ɲOaz�#gNm�;O��˘ť��� �&K�T��ԯ�lq�ZC��&��)T�}C#��)~(�oQ �z?����=��2�h1��e���	_�V[���?y>�`����dc����>�����k��JE�W�Q
	�ARU�f�(3���	�mz��y������'q��!~x��9Y3��M�@c���xA�S�mmEw�iӟ�a����l���<��]���EJM7�~��3�:I��t����*��6Ϊ�2���i�P�0Pe��"�Jl�z�B���v�6��#OV�˟���x�"`�: �1ov�9$�y�y5�T|��l�<\�^7\c��!�i�H�q�r2]�2,^�ڡ�P��l{𨌣�K���R9��I֒���9h/����zԕ;ԧ�a�d�N�_�M_���G'ᤱO`����<Ҏ,��ީ��
��Q����b{��(f�GS�-���,7sS�˯�9�����m�Q��(�$�^���ؼωܵ��VxS�T<
wy�a"\\�S�%��S�L"�?U��]���2t�����U�w�ꬒ���Ä۱#r_�Qױ��}��`�j���������o8L����I����/?GĉZ���^�#dP�0��O�T��j�D��s�w3�*6ֶm�2�(���R�gr�ŘU�\�Ñ��C��(�π��^����%_��ﹼ�<u�ߓZ�s�5���e����YV�0��/�g�`��CG!�(�^�փ׆|N_������S~#�>��)ơ�oơ�(�$�2�8?aO��0��sc���!n+*w�TȊu6��,�����x	��$�1브!�����]�X�윊M�S��ĥi�f�'�Y>�<K���|�F�}��Q�X3�;N���oѓ�5�/.q��3��^��e/K`�J2&$q��'e��&%tft��)�r3�R����qnNl�^p��sB�F��U���0^��1�І��wG��;�$�l�:Wy�"$��	�~�f�) �r˺D�n�?4{��)�H������xz��{�3��h:�g%�d ����d|'��"s�3;hpO"nM��}v�J�㜉W����q6�y��J:�b�>��<�*@�|�+��82%�g�|�"cLF��-��ei��3�K��or<�Sd�
j��Jڐ� _=q�%3��U`M��ʘ3I��Μ!�F�[�]	w7ѿ�+��k����Oo��<�/c����컔Wў�����Mp)M$x#
Y���U���y=��*�)�C{eP5�\�`�Z�qe�msT���ړ�j|�$�ۑ@Oi.SY��eAAiYv��,�����hr�ð����Π�d��sAp�s�ތ����z��rGVy�| ���חm����"�P�۲YL�C�#9 �M!�l�J�o�ץ}���<X��c�q��wbPct=�7X�!��Q�,(_�<<J�x)Jl%�h�_Lf�=Q��EV�I.���(�7>q���Q?K1�P�w�wm�I)���!X�'��V������!`h�'f$9n}W�Q`�2r�Z�������.���KvSf\����L��ǭ�<�n�|��1�S8dG�]j~��H����F�o�S`�\��SKBv�H�Q���:��@�2"�m}�7������f�o�k��`�{�@��0���(�MڛO�r�?^-�T ��_ʎd���&c�z��}�~����f@�j�(l>x�����0>�l��Ұ*�Xt��V��Sxr��:D08�#� y���(pG�x���I|�;�|� �`雔ӨV�kni�>�KX��zF0� Q/�%��#�gQ��D�^&Us�(r=�!��f�zc��H����^z�`����e�C`�<}J=�� r��ˀoI����Ճ��w�/�!P����Q[�Oun� ��e��6�rKX�.c���a.9�