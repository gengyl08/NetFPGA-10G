XlxV64EB    282d     cc0�P�� �W���At�@Ŋ99���ӟBJj������|�9]~:V�����M�8;X�%��`Ƕ��t�"�8-����@�X;
s~�dyͷ���<�F�r*$�o��+1Q��҇(m�M�<��{�Ĩg�g�_�!��\�uƦ�^�wy¬@���\�V[>D36ܒ"�|��?��z�M�<�˔���s�*��Eە"�`O:Fu�	Y��GЉ�/���3�P��c�������6��i�L�mf'.��`��P�^.&f��ՙ����
�+,���}W�3��+�� _v�[��q>�����>~�#���e&�ΰ�:�$�b�y�����~��J'�OqWO��.(��#�7��~ʏyTNW� s��y�?5�Uo��1!�#��s��[��_������%'��0���o����AY��.Ҕ�F�0�і3�G�)�����l�����IP�W
2EjDpye� q�<nA�d���o]7��c�[D��M0�*S[��G�	(c�9�o����$�t���P�Ʃ BF佯�	KCh[}���:)$��{O���k�1#@ˀ��]�8<�^��|��]��pʟB�x�`���1�D��؄1��'�Fc�p�=�m�g��m�rMKS�>�y\ۏ�{�
��x�d�ȫ�����D�[j���Kj�.��#�j��"��]c�kcP]|�)CX��ŭT�@]h��1����:
v�Ov��9����j�A��Uي�yc�{��$�wı��I���6o��ab>��x ��l_�SP�ܱ�/"㰪0NS%��҂M[^�Yo����p�9j@YrB-Q�9W^ ������u��P`Zi���Wn)5�xl0qw������f,r�p�){��@|:v�1`E�b��"�$A�8�XV���{�r�<ȱ�ғ�l�ZH/XC�#�P9�#в�5���j�&@�V���Kϼ��C|����}=-J�t�杋�䉅@�mO(`��O��1�	<l<���6	\;�I���b\g:� *4�� �i��˫���M������=/�G�=�[/բ�}��W��:�
ϊ@á���;_�f�M�4�=Q8_c���	�>���]\I,v���G��c!��l1�́^��X{d��7! ���\�a���̀C��*�il���?�E��
U2z1��F����?��*��P*�J�Q���YB1v���k�k�R��b2�����ǭ�D��n�(�F�����3K0
A[>�:1��2��E�܅�g�L���C�M����$A�7���i���wE�Z�����3*�g`K��~�R\�����:{Pׯ����9�Y3h�$W�I�##Mm_A�}��=:����ׁ^�o����ӗp�3����tki!:�x���4�j�`�g��T�������S_z���$�!Z|�1<fF��8̶;����Y�p3��G_L�3��һ������u��S�{�-X����/�{׏)΢u����	�v �K��ӓ8$��S�KR��Mp3|��B[+e#�uY-��vWr)'�C�O�,���x�'��m��#1��k3xM��-7��U�u������AL�I��+T���Pv�E���W�ŀ�f<d��Le��ˆ�9����U�WКgxE�tED[��#�iR�;���<�q~t�I\�Vɟ=����vXE�.�u�hV���r��jtkׇX���p�o(���{-��IS{4Ck�$�:��:���B\{����0���p0��������I�����O1�&M��,ì�����^M��8��K�A.�q�V�bj�!��#Y�^Z��䤝�\b�$B=�g�����d��3��Hv|��c/��v˨�o_M�p4��ܰ05��3�Lb��E�G߳2�l��3�4^��Z���7|:�S&(f�پ6����ў�>$���/?�v:ñK���&�?Nb��z�cBNNENa'B�/���=�Ē�iR!=����J�F�f;*��s��"��`�G3���I�z�o3�КZ��p������YF4��@EJIn��>m��p���İ'd�*�G��ᒸMF�=�*k����b~�|dO(X1�t�[�K{p+��iP�#��{�Wr�տ�_dA��w��_țA�^H��|��՟�ӄ�y<,���	 ����]�15���;�Y�����Q�p"(x�7j&������������娥¢�{Қgtw+�7���_�h{��QU<:^�.�t߻��#�m���IHc{�R�U
�i��e٘Sa%f�fc'F��ԍ�, �Z�����(|5��ic��h*X�%�y�+��(��U��p1x ��<�)^�1�uR�Y��$b6��a;�a
d��B�K�*�ͳb�Ȑl!2�����bE���6���O�~���>*��_�]���<��[�d)�_#��%�N�q("���!�:�[Im:�jl�^�{�-���sC�Y� �G�P�8�/����h�8(!���x$�rA�ԟc�a�r8��:)�Y���� �=z�6�ᓥho�(J��Ӥ�<sp�"��L'���:�TY4�Ppb!��Ul�y�/�)�q"KQڶ��1�|�|bf�C���T�=QWX���D�&�����! 8�-D�p���QƔh�(�R����xA�W���8�M�A���Wt�I+�x�?�I�b��B�њ\I7�B�z�Y�;�$l��������ƛ�<[�ov/�!\��.���)\�eh�qp�H���7�~\�d�) 9C?w�)E�-�!|ć�>=�x���m�y�)��� ;��H��^!N���Ӵ�zmx5��Ar�3�|%�^�"#?���7�r~�z�����i�҄|T� 	]0����J�tl�z������f@(��08ctz��8l�h���s�|QR0>H+��㌩�'4��v�ܦ̅�^R�|�pB���p����}yR x�v��Pz\��%�5y&4�[�~��J4\~Q��)��%�8/aJb�F�_c��nN8�uK����������:�$�������,q]��{��R����zG0�&l���5&�eB�u1�٬�N�3�]A��8:���s|�I`h�܃�8`�R�_�?Չ���� ���b`�O��1�ݻr����ȗ@��0���`'��|����YM������avq}>�������M��"=�26�A�p8�53��~���[fS^fA�&�
��r��