XlxV64EB    8a6f    1520V2z�|V�.+���#��Y�G@���hR[�E���<>o��H� �u� U�� '��c�ڬ��,���OK����k��S��;��}]�JUS|��-=k+������*«�(ҏ�_��&�jo/�q����oF��7���["�r��@���q�O��C�o"�_�����'��%f�6Q]�J�1b�% Γ�K��D�e����2�X�a�}��&�yN;�dݬ����<$�î�����r.�,ib%t��u�&~b�D���L�SޢA_��Q-���樯������}K�Ef~PP�6���!Y�����rC�G��]F���$qw�R��N�[�g�WPY}ޅ��Vm�j���Ƿ*Sٹ�)z�eܩr�`&'-p�?�$�^t�+0�2?ӥYObp�o}� ��@�|��J�ֻ�w��Ben uV��I�����$T�I��S��9��Ct0�M��c�r!���k�w�uIl�).pj����}p�$���br�V���Ր�<�l����9\���1� ��6�Q?-�����~�Z��utFȒ1mO��\[�����?F�.w�i��c�$�6�g���n�;/:�cr����?
*�ö�W$�n���P	2K�Z+V��(�"��u�V�h��-�<�v����'�4;�-ҥ����E���A�#�;"�$4�f�C7���Q���ou6$m^pN�Ց���[�T�p�n�+ ��MO8����hAСQ��^	���W�o���Ӎɀ�˜#P{�q�o���
����C�K*@�H�8�*�6.|�2ez�"��|B��nA�Yϑx%L��r1["r�>�Օ�W;�9�~3��Ke%r�l6Ivz񥾑��U~�~R�6��p��c��k�l�p����h��\YԦp�s�����^�nF�8cjp�k�W�'pL'+W�쉛� ޓ>�ڻ��2S3���3�LM9����fF0dX-�k_Yj�;]Z�<�t��v7��uA5vkٮ ϯu4��~�K��?� C%���ُ��Z�t��7�g��b��d�t���0�m��x�`���9�D��k���{^�����Uc�����8s��c��HI��?j�W�����n�������q�O�i�Yh�[
�g	 �e��-:��H7
��"��A|7ļ��a�5�V��-�7�U86� 
Mf&�rl���>GW�85!+u�3C�~N�{ �<��n��exvyl��������m�	d���i��c����B+]j����c�HvO1XIG.c:����t0�x�5�Ёd��u���Qȁk��t/_h�*��*�}Y��-�,��Z�E	el%.O�2)&��:�Y��~�+X��=`�]'�O��ޘ4��XH��/x��Uq�
�dQ��L!D�5O�����bi�:����-���y	�6���_K��J��+�I�˚�7j�%�}�Lݱ�:���ìE�&��Oh�X؈�2������qhT�ϝ����xgvB8p#x2��˱�(�>͕�(cG��ȵ%��L%�$Tf�:g@��s�e�W2Ќa��X�A?��'9dA�zӣ�}-@a��(*Ҹ�0ݼ(����ݬ�0*Le��-3*�p%��G��C��VyE�#�@-�����Dv�����'T�����z�}�2+��gC��r�v�,�����=%��u1�J�2�7�]�@�]l��JҰ���[�uI>aaq�������?�����Zs|�	T�p�wz�Ys-�vD���{C^� 7�����U�.@�}yZ_o)�v+��t(�BtP��E��O�n��\_��+Gf(�{��D��M�e%�4�lٹ΋��4�t�Ѹ�pi��U�d�tƮ�T����N��-��7��=�פ����piܵN[C��[�rQ�ۺ)��fs�o`ޗ'5��_���꒜ypr6Cf�W��}e��l�J�s����w3"�bW-���LYEV��T7*1 �nQŀ���+P����Gs��V��~�v��5m�[C!���� �D���5͢9.��՝\�!wM�^�����.�j\�v�I?z�f�ܷ��	�?^SH:��D/;���KBR����l��@�yJ6Q}9pY�I���vk���{��)��`&���t|�p�����.�	6TJbsT�K����K��rXP^!X�����zLt�p�{Z�T�SJ/��:��	�	���b��e�և��.At�b�ӕ�x���Q�dBC���!�Wtڮ���9�A�sVmSw�!#�O�D�������_ ��|ĵA���G� +C����*]���!/�
;�cF�>1�ҝ�}0b�-u���fM�ޖV�H�3��3�2�i8�s�ׅ[��|fe���j���f�:���#�Z�XEH@.�9|��8�{O�إ$��8z���A2��J)T���\���ޯ��c����֤��D`\��EX�,��������L��kT9���,����V0�4������4
�Xb�W��!��E����Eђ��^�<�������5�+����h	���m���.T���>��zU#�(�{��G#�u�3�z����~��Q���S�(�c�j
���sSCxx[i,(�~E3[H�y�<?�`���}����v����qi����؜Za;��6�+�u��.
O�Q���]ʌ�w�g�%�����~<fd�ʭ���:<��k�7^a5[,�zz�J��*��}���uE���dq�l7��ۙ���%��5����{s�0�$ff����TB�����jɆ����%�4�9OxA��� ,l��T �<)�X�T�ٵ�L�l@'��:���
$"�@K�~���aﵞzGb�S���>��x#�����£��'��>2<C�0=R�U��[�[��wP���	 �j�/� ���	üӇ����r)�����]]�Em���,�\U���4NN�p�:~�(]����}�RhnC�y��U6�W����8�{���uM�AB�+��P����8�J`�T�:��|��7��C��%��麚W.+A�-|N�NT��
(a O���Ile�艘�����ł	@�~�ڍTn���,���|V��g΃�_ ��qd���@A�%LNTJ�*+.�?�lF��K�Z�<i^�>�A���8S�(?*�}n%eDZ���mX�z��J.W����z���� p�ߪ�(�-�0�&�J0E1�[�h����Z�W  ���!Ɏ�9�}���!���ՃH��=��;,Tzβ$�<Q�x��=l��VJ�*h"�R���P�}�}:�� ��'$0!�������07��]�g��[KꓶK�̏4"����FC#`��y��}��7Ғoyـ�f�ʿS�~�\.Ջ�4�.�����r���{��+�Čjk�Ya1,����Nb�F	��n^���z+�gL�0Sb��,��"�8�f־�R"�h!K�pcI<M��SƆ���H����YNI0G�vy��rA�*�¸�d��/���xf�mא��,<$#��M�'�Ka�h��%_A	ccN�� ���N{/�N��_m��=�֪��?�r�䒧J�-`Ш'3�造�a�S
�{��]��ܒ{)��4sK�2+�Y#�իg�l��)�8]���
�����o^���w+B.���`�hV���� ���-�/�_�^<[���m��"Q�2����!X���琮�����F���sE0�m���TL8MXj��������kN~tne}��%m�YJ�&�Zs��qR� i�5
�=�	�fb�B��x|��450g"1�q.��@g�׸�99@��=�}��C���L�u�n�Du��LE16��S�����Q�mjNQN���.\����������{��0�#��7�6��g��֢�+�Sh�4�:(z��!OՓ���3��ܐP��9�8R'�.�ӺN2G�A�R]�JW?F�E��59���a�UA�%��v���-ä噙�ȓ1�S�N��^ �PI���,N��h�49ϭ�>��׮⠭�����?b"���~����oYճ�R�~D��}D�`m�$$��E�'�²#A��#��'P��w��RI��gE
��`�x=@�G ԯ��GX�t�N�I1.�V���	g�����+F��<6��  ?�ޮ&�ﳨ��fw��YJB��n�ռ�2���Ȓ{	F�E��mO�k�L�<]d����=��gf�A4�aUR⌘���UjP!b���0͜�.�ʈ��4�llKO��s��E#�-���%�G>��F��m����*3e�XG�mj.�]�����O��eנV�*��4B�ޙ� �\!K�I^3t5�_ⴭ�vf��('��6;'��Ss7�YUv��|�P�(�N}�bOH�P)����(Τ��]�� o0A��o�o���բ�E(O�7���ֵ�:"Cgn}I���������.,����g��{Ű5��%��"�In���8Sʉ��TM��\�W���[V�~�!�<�}]I~��z7�TA�Cx��	&Ԝ�d����g�o1ݱ'i�"�ڑNO8�]H9
&�a=ox��j�3Bꦷ�q�O�Ca	���Q`É����u��b0��F������l#p���A[�6��(�޻��ץ�x�1�C��㭜�Ix�r�v�f�u������ml�1V�������,aL?/�e�l�\_�ɩZ��}ȇ̚�4��e�:��P�����f�f�CFĨ�y#�@�bXg��q�d9+2�S�]��y-$�ޛt�1T#�5�s�
b2���t��Ӫ"�h25��h��ZM���.�:��֩#$�u�|�'4��)�eH��#������d�6��Tveٲ����VD�a%�,%�34���L֌�Ge��5[�{��=��|ɒ�p�xgɱ�&6cU�'�t��Ik�sWG�o��{x�ן�6^�v!��q���<�Vm��9p�뇰������X�h�|C$�
����ؕ'e�fU��6 ����l�U���:,t.�+B�tFG0���z��m�����o��EoD%�cE�Z�����D^y��y�t=�s��d��V;�D:��pn|�	������c���Jܐ{�E-_]�Jd8�t�&vb�Jİ���b�o��֒�Mf�!Ehi�r+l]u]�<�(�P$	T���ux�3[0�z�rGOp?����u����{`��^���r�ޛ[Q��Z}#��wb�������]n��)��������������f&b����-�E��Kɍ��]F���%�_Ynu�KT'�1�|���^������C$Sb��Ϧ���%=C��\C�}| �� k���M=��r r�˥3�k�I�>�� �DI�;}!PD<�O	'q�_䔼�͜ƣ=P2�)}��%�ui�K�;�V�]	NtnI�x�#@��s