XlxV64EB    15ba     850�N6��8,S�+�U%�'�Vyp�����
/'�2Ƿ�}*#k� [p������S�A���5����5�=���b]������0��h4A��>.NwTƭK�h�(F�p�*��M��L�Nk%����P�SdY���T�Aܱ�..�>Qq^�'xs���K�!{�`�n�����8��<���@�o�����t[���̉6�Wd(܇���[�����z�]�Ү'�k8.-b&-��~��s�cM��1�0?	W��C���.�����xž�v6��A�p���?nj\�b� G�{}!����8�����>�4��P->�_￞n��-����9Ќ����$��ۮj�X�A5��nK_��T�5w�b��7�{6?��3xC�e��e�LC�vWn���������l���aS|w�3�=܆������r��He���į�k+%���W,���?����%G��X������}%��7�,�r���6Cgשc!���0dWс���ӢF=H�c�����r>���q�m����k�ٮ�[f��ц�Y���[�b���k���1������POTq?.�P���z˭�X�-��V�mW:ݴfN�� /�B���Ԧ*u.�Za�$�(r�9�������p�j�v�1��F�`^p�z�8���C�� �X6Z��=�j�H):����VV>AϪ&���du"XΡ�p��M|�j��5/8F���X=���[���]���.�n��l�n���+G_�Sq70���]*���;�*���h��fOb�o�8�`9�YB��BZ��l�/i�"�!�[����Q�,*�>_��A����EJ���rY]��[��b9mX<�f I�^���=2��Ȩ��Lp1�ت���<B�U�:�N�=�MgM���Q��8f�Q=���V�V����&ɞ# H�-�h�a���g�'�ci��@~�\��^��DmG4����MD&��~P�v᝟9}�,q�8d��i����Lh��uݧ��2*t�7�c�I ���m�!+��ڣ��ͮ��X&�*�OUe�Q b�豍�hGi������0w"�?�3vvE�6<2p�[�^��ˊQp@y$+>P�� ��k�k�&s�U�e��N��<"��-���]�+ǥ�~Q���(�,����x�r��NQpD�ɧL�务�P����(�@9k�5L2fK��Y�j��g�7nP�,����ª%^��y���>����E�۸δ�~��i�o�#�l����:TB���?�2�����ϖF|�2�wҢn/y�� K>]��_\,��~	�x��9�9r��n��馜����C�U����ͤ�P��^�X5-X,�n���e�;]�Si�J1 s�_o�K�lY����>����pk�~Ͼ�pL���P���
(p���3�n捩w�Y�s�H &A���m.��]-�<<Œ�D���ڴ{xwy�����%Ǫ���.x�-���8}�����p΢�����>I���E�Wk�Y1��PSϗ��ya>�d)�5������{��wdJD��]E\ˏW�Vi;�-�}����k�[+~�:Z��/hI
�e��~�Q��|b����a��j�缸,J���`�k{� Ψ��|&	|Ӏ�(�����Gh�D_n���b�_�)8 ���C�E� -5e�ʣ���S&�G^��IaI�����O���}\Z��;�C:Ոar~� R�hy����K>B��@I���h��3B�$vn�N��x�����ǉ�E��� �.��D�^�$T�q�;)�����m+�/�䊗��{w�5���� ���"��1��
#n��z:�'@�j���@�R�#�s��՜7�����
Թ�j.��!Ñ�|H(��y�絽	���1���&ǵ߆���z�j�~��UF���0�`m��HHa���sb��7�i��m_�a1�/�N����=wy�ͥAH���Z=�VDMzCVϛc�]���!=wMx���z�=Z��?�e��}ܸ"d�tx� -��qN����@j�w�y��#�s0K������4EƏO��+ޏ�γ��Nt��E�����3$���FPe'�