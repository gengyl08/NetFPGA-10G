XlxV64EB    820a    1460C��+c��̝'/<S�ߑy�|�c���	�G�R��L�I	�tw~���$�x|i����
P �`H�y2�vY�Ƥ��qI���B��hO>N�s��%��Մ�Ÿj�&p��'�Q��r�|� ��!�B�E/C�:�ܘA9��'>3�Kx��2�p7�%��ّVQцh(�FFJ ɗu(�m �=!�1g��v���&�|c�h2���l�����}�KEAz�Cv�B��E=f�;9�u�#�.*��liQDSL2�n4�R��#�a3�`_	}&NΎ��1>��c���N�d[o�xlr�o�j�jY�P��0�H�O��1���0e���&� ��Q��Φ��\��xJEЭ|II'����b��������z�S_���n��h�8���9���e�@�n�w���y���|�&C�lh��h�!D���r[]�� Q�L�$��)���5�2,�,$����[��$/��c�T	���#x�R^��{?�A<��2/��4[�/���>�6��3�3�j��:�5�+	�Zг��b���p���uL�B�&�q&��H�yq����~�=���	\?�������׽,8\���u��tAfp�i���4���a��s�-2*-;Ӵtr;}�N��cZF:L����ߕ�ƤNM6��R��c�z/B�0/֛Al����h?.��y]J�g ��:N�QP��i���P � *��CK��IL��S������{9(Vq8U�ǚh7�\d�?��2�tK� �
��Z(��e�BZ�����-�T�mO���8��c"�������U�@1�N��:��(��_�0�Z^Pn�rs!߭����O��Y\E���29�\��4!r(S�%�d�W�䧨AR��N�OȐب5�@Pk0f2�2\�3� ?O1��X ��*ٙt�n�-�~f���}�;.]���XI��Q�tgP��
,vg��y��	,�=����.����lP�o�#kw�%slHV��#cc!k���"�l6Q���w!�Ir&�d2@c���%a���n�)W$����;!W���^(��g��dp��3B}�]���g@�:Tz�L����s+}>��`�5�虇��O�w,�ʧk��nmr��?_��S��2s ��^����<�����v��K��yz+{n¼U^�Soh}�Rܞc���09��[ڷ���������@���r��`��cĶ@��5���_��Q�=����}�6�.���$�AKuk��+)u�gR!8"bY��.D��sǶ�O��V1߯c\=�j�v`N�9O.g��� �It�uҼU�J��1*� �T1�s�cT�CE<?�g/�-BF���xN�-8&b���<���E��~���٢N;9/��8�3o��
��Nwr{�W��w@��3��(+ u�+�lLG�G�0�^��=�ӥ��'�	�����^�m��yt�� h���02D+��&�	L���``�����KE�CT�ҩg��Ow���������/��et�1:���Ji\t7?��)�^Йao�3#�]�X@<�1I~��.~���W
��B= �T-}m�^�P���j��.W�b�$��D+�i��C�s.�X}�ɋPb�d��_�g�*S�+�m�P"H��jf�G��9r����cV�<&O�9�1k#p��9���#͔�|�
L!�ü��#��i�������m��hy�������L�`�� �գ<����=1��KQ���1�l��d����[B��T����>6J ;�S�>^�҈���"{	KJxg���((���`\x,u���e�R�r�p�U��l~�1�+���R�%:*�G��*�{?O^4�ol�*Q1s�͑6/�X}d�ȗ�P�Vs�zT������ޓ�]a/Ή��5}~��v�a��e��~����0cd᥵�z�ca��y�^|e?ss�/gQ�\VF��)��a�����~��W�y]�6�s��w'�`��ް�_�\e���la�Ɯ��.\�n��]�u��Kĳ`-zu}VE8�iTܹs��'�05e����:��
�!�a2T�B�V��Y��N��E�_���1�8��<�!�ʑ�o�ɘC����Q��-�$ۮ0f�W� �<�o�\�0G=D��H:��:�>}��N��×�8���g�#��R��Rg�_�c��7;��?�7�� 8m�l>�V��5�Y6���P�[�赎��h�6(��SUlABԼ�V���mdWπ�F��=�{(��ʝh��x���XG��/���*�	p�~��
�&(F��B%=y��Rӎ6��?��׋R��y�[�ӳ8֤F�o7�m&y6��H���x@�����Ev̅�f+��-�4�a����$t!�E�v��2�TT������n��a`��^w��.����F�������&��E���ߛ�J|���VW	�o�����ܤ �ٵ�KXkZ���g�r%5�I9~L�����z����+�$JI�)�KOM���`[4�ǲ�h+,�U�16�_�	[�D6U������H��'��12+�@�)!��2
��Wv���#y�;%��sq�.�4�Ӽ�\�!H����:?>W�/0Taf�ȇ�D	�:n;s�z��?,�Q��El1���X!�ư0��r�DU��+���ς�wRr�R��MJ����s�!l.4Ӹ&����VRC�!��JF��a�R��B���B�;-�?���i~L��ʦse�BL�bA;gK+9�V�IX胪��E��3���H�.���C�BC��S{a��Va|n�,Qg>^��T�z4!s]���0�����B��@-F���-��e��m�$ˆ.��߂��5[}x����yͷ��e�HO>\1xr ��%��.v�?*��#�+Ha�<6_Yq�J��O����#�l�դ���Ep�����"� �I7z�&{�?�k_�
 ���tr���&�ļ������� � ��0���\J��Ү8��7��»��lx��ߐM����D�;E荱�2Y�	]�3��`���a?�s��B�������Q�~K�Q�$a.�c���8eCX=_S<{�kq�����rA�6U��	��OX�����~�҅���zS�0��CoB3�1�-П��V!v��g�l;Y�oND׿ߧ! �b�
���ijU5A/�ݝ%-��wq�C��Sf�^���Ymn�b�-/��D㚕r���sa�&I� ���A�/?��vE(:i���O�`u����<"�lu7`��b��W��|�@i���ل0U�|����ٞY��Qd�ՙ��P�\�O�w,�(,�:ў�&��؋`n�SI�,#����
G�ڷ؍#;Ku�zO{T;�^R.�jP�-��C�qdT�ӳcn��dGVn,Nz��3|�̅=մ��	��_���3	O�9�d(GT���.IE���L��ȳ�:3�!;	,�W�d�I�_�Nϕ�]n>V������q\��c��=0LՂ��tq�'-���lk�p�;x�dɄ7(U�jש�&���)��f��?�}���s��}[COm�(H!�ظo�s��7t����ƛ���i� �n�{�,|�	���|��gd]�U~=F��(��k���Z'�]_�y�?��-�,�Y ���y��T=W/8�������{(�zH�Y�RShv�g�O��F"����0�U8��s��n�M�B]�c?���8��"�r���2�G+R�Sh�[������*���u�c�T�F�˒V	ߩ{�</w�g^Z��X��n��@x�49)M�i��e�d�
��cw��w?8� |r��h�d㵈��p*� W/o��A�@>$�}ǆv�K�G��=�RfE�1�>��P��T����Æ_���j���+�F��Ac~���X/��V��@��
�Ph[���ߕ㢎2PR;�ϋ�i��Ў� ��L�z�K�:����I>���v0�(�o�w���e�!��<�d�[E�r3��'hL�0�DJͨ�9�K�NB���d�H]�Ѓ#N-���ϴ�����K�|>���9cێ >�l���+�QuL{s�)�[
>�kjǻl���/rYL��nw��b,P��H�kS�<���d��x8��B��}4�S)�ߺx��}B���t
C�$��0�&����3��<b�]t?�0>;�~Е~��5H��C�>������ĝ���M����29����!��e����+Ɩ��%5�����o�o_� �*<��s4:(���w�m���)��h���I��h���U�zI0f��l�v;3����/�K�am�{�V1~��%�6�4��OnvH>Ќ�A:�G�y�h[A��m�L�����f�]YLȽ��CƐ�s���n_0�䜨?��7��V�͖�Cy�� B`����J���?��x�=�]ٟ\�G�e�$�]��A&���O"��+$앆0�Z����>"6���ɲL�)X�F�e�^�R��J���s_���Z�k�X$�t�A�!��;���qY��V�������YG%�uס�ͽn0N�;�	/�N���{�3�fꢅ����I��b�ȩ�5�� �XrN�a�[,�(W<��zṤc��5^1}�
^o����kalX� ��;�Kl�y�����m���"܌N)�畼�e+wXz��n���4z�?�� ^�ƙ��#�AK$�uE:�Z���{�L���X��Z��'6�L)��6~
�f����P�ZJQ�ʶ�%�R�2P�
��� Y3I�m �4��<��� ��ym��yi�|1��}��t���(�Xع=�6<�ɭ��ϒ��#i��\�7�;�H��l�� w�z��y��h��i-��½Uk�t{`������R�EQY�,�ۡ���Py9&�/�9 �ܳ���I���	�FË&�L��taF�#�iRwJ���.�ɡ�&�ߑ؉Bc�]!��Y�*}ˑ)'\~`��+�-���ܯ�$9�LV4��5�QϚ1��t�d� ߺ�nG�u-��0�-~��P��M�����z%�t�4#L�=�x&p�s����B۰;���t�$�����K�{iUj��c�^����9�P�!W�(���a�`V�|��ף)m�lKYX���U���