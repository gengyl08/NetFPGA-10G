/*******************************************************************************
 *
 *  NetFPGA-10G http://www.netfpga.org
 *
 *  File:
 *        rld_defs.vh
 *
 *  Library:
 *        
 *
 *  Module:
 *        
 *
 *  Author:
 *        Muhammad Shahbaz
 *
 *  Description:
 *        nf10 rldram controller
 *
 *  Copyright notice:
 *        Copyright (C) 2010, 2011 The Board of Trustees of The Leland Stanford
 *                                 Junior University
 *
 *  Licence:
 *        This file is part of the NetFPGA 10G development base package.
 *
 *        This file is free code: you can redistribute it and/or modify it under
 *        the terms of the GNU Lesser General Public License version 2.1 as
 *        published by the Free Software Foundation.
 *
 *        This package is distributed in the hope that it will be useful, but
 *        WITHOUT ANY WARRANTY; without even the implied warranty of
 *        MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the GNU
 *        Lesser General Public License for more details.
 *
 *        You should have received a copy of the GNU Lesser General Public
 *        License along with the NetFPGA source package.  If not, see
 *        http://www.gnu.org/licenses/.
 *
 *        This module was developed by SRI International and the University of
 *        Cambridge Computer Laboratory under DARPA/AFRL contract (FA8750-11-C-0249)
 *        ("MRC2"), as part of the DARPA MRC research programme.
 *
 *        This module was developed by SRI International and the University of
 *        Cambridge Computer Laboratory under DARPA/AFRL contract (FA8750-11-C-0249)
 *        ("MRC2"), as part of the DARPA MRC research programme.
 *
 */

`define NF10

//`define EN_TESTBENCH
//`ifdef EN_TESTBENCH
//	`define DEBUG
//`endif
