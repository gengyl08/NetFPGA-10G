XlxV64EB    431e    10b0�e�Rب��r7�Y�bq^vx�N�p5'ǹ�ڳ��7?���ɜU�|e\��@�����ZA;S\F�Ԡ�6���=�C+T��c{�?�p&�ٙrM���-�ї���������!2=z�&EIJ)A���b��o0g9����7�m|͞��ѯ9�.ݍ���WR���P��e�TI��'�A��ʝ�wM�AM:m��ssЇ�X�%�^���Gu������670oH�%�ꒇڡ?�_��.{8P��kz�LD�<�x64��L���į��?3��b�O�pNט��~�\���U��������z?��3�4�aZ^t?2-�����$C�t�CAiP���D��R\��x���@��z�N���oʐ�)5}9��j�iWT�e�3W�I�yxD��"3	5n�X8iU��Y6.�b����D��[�ܤ����/��}����V>��������.XpEF����^z���M'"ޛ0���
�p��ȟ�1,�*rG�]���~��-s����O��/���PZ��C֖�J�r�*�+9��4"Z�ҿ�fE �/ [�Ȃ�7	����+D��JVOC�^=6])P,1=�z��v���@�f�&d-�ES%���oR�>�)CL���b��g�����?ܔau@��T\��5iŷ��Z��y��C�<[s���3B�A�-��z��-���?I�c�?0E�DnV$V�#��jZ����!Q��B!VZr��ܴJO���
=���iAF��� J���RG��3�s���V�!r̛��3�j��R��V$�l��� 9^o<E.EZBs��(U5{`�� ��pB�x}�~{l�2��bA�<��,�Q#�R��/{^����r�����5[����hB��� ˑ�"�㹜ۘ&��0�L���z��.��R�A��^0wc��+��9[��lvT΀ �F�E�ި4Ղ	b�9@�x�� ��@��'�X�����.���vܩ�����dM5L��a�[���6�>O����6��,oyI���4�i;Y;_�0֢^y5��-�����t�����
		��ݴp(t�S{0���|�"����egȡҐ#������'=��Ϳs��6:"���v���RwZe���R�o9�i���v�DpYbA��*	��m!�H���w�_z5������r�i���lޱ�=�yj|�*B��8�y�j]��K�fL{3�msɥ�Q$�nѶ�iMR���T!|ŴC����j񂋃�x�<�ɭ�>9zq�MM����U��Hy62�ޑ�[���F���t%��-�)«�G��4y��l) �ͪ��P�����(/����-�Q�Ѵ�{��ܷ�:�H/�����t$g�\���R��z�����h��O+�A�����r���U�/ir@3�R[7�~c�,�M��Gm�d��u���]�)���Dh�JY�t��dj7~O���X{�-�;�KS$���u%�׆M	�'���^��G6�s�:~l���'w��຤8Y�@����_�x�VC�ɀ�"֑���6Fg����f}����5��Z2���,W:��]�F��txk��($]kĄ&�=vJWt����թ/*�F�J�UE��V��F�/ܫ���j�Z�&	�Ɇ�5������^��jE���N'���}�_��1�jd����`J�%-p�W��� t��晽^ŕ�`z�[S��T�E���k$PE�1\5�pQ��8�ܸ�X�����#�S(�ג��%nI!
>N��qP����B�h��R,G�F���@��R'��.͹_��R�$E����	L����<���'u��:&�;��*��~oV����0�Ы�x
��z�=��X����"���Ѹʈg�D��T8�i�Ɔ%>�s�� ��]���^/�h��
]�.�O�H8��Ε\����b ,�1���	3anhR�e2]X;��y���������F�f'���Wqw�t�����Ze+zp�e�{ʠT�^�\��]�U�K9i��y�C�{{�e�����^v9��V	���;�qm+�z@�]^٪��ʝ�#S�&`�J��B����Ԙ5���_�1ew}�C���:��X�u� �V�h���j)M��kZK�N�M�"c�R�6�˜LNvڃ�󜘫p6Ź�����:���`�J�n�i1|�,6Ԅ��~�O�R��?IXq�w���D���ߧ"�8ߋ���Qm�ǆ^&�G�x��|�ld滳����<;�o�7��}��3lm�ݭN�^�>�;��X��Q�����e�x5�<�����(�4��N�~�O����'R���R�S-%y3�*,�4(WR,{��j�'a��Q�|	i<�{"G��0��JVr�
��F��8���3�ǼWX�]6��x��~]`��lM�ͧI��ȝ�i͂mdQ ;�n�8���;Q�%�8�!�Z��iA:e��a��i��"��;�
%�74�!���흉�;����BN[RҚ��{gU��'���K���2��"&#��k%o���.��P��`5��)�'m�M){xL@�\�� ���b`�%�{a�k#�\�oU{�ջ�W,���[�u/U����|����S��k_��I�M��c]��[�'��F]�Y��M���5��tIg��1��d;��6*�IuG�s_����]����nE�>��J�Ai�	s��'FL�k�A��_M�Њ���d���;܈Z�*��D<o��6�w;�+�`�7|��҃�g���uP�P*XJԽ�ă�Vp��/�'��6������$�m�@�C��ɀ��^+uӬ!������	g�o)���Bp<�vȆ�T�4�Fi(�~��W0��G�>�Ţ�����<�^��-Rd )�B�G�_�����:d��\\&�7�P2x=@ʳ�Nj)�_!��$bf�H@Et���у�$|�̺���Ox���]��a�6G�j��4�i/��Z�&�L9��^"pM�%�TE19�TO�\�{pH����:U?'�j��g�{�ks��
� ,*�c�����wՅ�����!�ܕ�F�:�t̨b��훴H.@���t/�-�&R�):�A�^Y����V�
H���zvQ0�
� "�ZϟǔOy�r��[!���|%'���K�m��7�$����tL����$#�Ǹsd�@�@)����ns�]�ͅT;]�6�7v��sU\N��=;0�Tc/	�������j��܆/Xě�h�W���4�s�:������Fy�4����j^;z��C��q_e�Mi^����W'��6:D�M�<lv.�g��Put�����r����)78���$���]��t.?!縍*�ĥ3M���J=>$'�W�<���|�PZ=y��y�D�b�����@8�}��|�-��/�^q�:�o]+�M0Z�H���ew�$���}�a��s��}^���lk4���V���=�3h��ev��7��=Q�a�'W�u�{�p"��[�ۿI�:m�7s��Y�H�^�)�{P�ȗ���g��,5�}:b/(�X�7�z/��!g��_G6&�\O��=4���wT=��=X����P.ߙ��Xo������ͥ�X۠X���I.7�):�[��U�NV�~���Q�0��g��M������>q��X�?����Dc�R޾����e���u��]� ��*�/�4����ML�.u�Jqg��f���S�Ϋ?���a�v'����\���>�d)��J��{p����Ւ��N!�SrJZ���>v��*����]��ғ����}��x$��[�]�%�X�����"2�(�ً��L���ֿ~�9��¡��ѷ"GL�o\��_m`�S tMTBҝ��S5/��l�($G
c��i�B���7�� �/��1��(���ꮏ7\��#�#�*���☾��eYOWpm$	�/���7������2Z�0�Ə9�SGϋ�o�?�0��"K��"��ь����;�k��cAq�{ɺFb�wHS/��j���RKa,���)�J�rT�Wg�6G;0��xV�!א��P��d�^�n���/�p�-�������fo��
ۄw�6���$�6���`r��dQ�s6r���OJ��/�d�>����Ktqld`�kl��QY�'�T<#{�����NIV�A�M 뫒��m��ٟ:���J���%2��u]9��%���#��)�5���ߍz�����.��#�W�&STG����h(��K�Qq�F7AnH�