XlxV64EB    576a    1430��Z[�v����h0.B��E3���*4\�Z�Y_\o���٤�@�z�/��e��� �i��u�����:�[	��]�&���q�<s�g�N���>&zM� U�9L5OaGFn�M8S =W[����b�5/�X�|����Z
�����$2b����:�� aq@KS������ִ������r��к�k�����Wu�-�1�V4��9�ځJWU\;���y���T�U=�A�
�ø0����G��05�	��AI�D�����j����^�ͯ�u�}��,T�B�ԗ��j��\�K�c����c6��j��9^�!��#꺂��]e�%�{N9XvI$�
��N�cP#郄�L�m������C�Ց��8��EŜ�H���8��{�9aDPWD�sk` =P`�a�MjX�T�TZ��!r��ƥ�y��%���Ｋ$��Ï�~����Nl!ET���RG?��wv��!���+^Y�L@�\�����n�s��x@j��ʀX��Ij(R_�g��A����*Ȋ!�/�M&�붳e�,�;g|ӄȰ��&����ʃ����7�/ތg�Y�S�kS�V�R���ЀJ��]TJ����}���]Ț���Ď
܂�;�w����(H�@�-�QF���b$�7�ЗRѽ�9��r�w=�3�u�&��_�h8~W!:?zS䵶|C�0M�ʶ�J��B&;]L0�W���,P�y��G���KY���-�����І/��i}�����;�U�	�]��E0�1ar��R�^�����@uƕ�X��F[ϸ׻�ɀ��G�/̛����
 4c!��^��1��ai�Ni�amO�����n{�c��5U-\�
�	X����^����r�~�w�d��>x�7�DCL �}v����W��ܚgھ=(��߱��f��[
�[�^C>[�峾ĚHc[��m߄�����,�L��bnP�Qϖ� TD��0�������Ol3�3�W'𥡿<lfLˍ�`����Zx����R��f{C��l�`Vd_�K+Q�BC�d�o�|�l׺2�E�w��ŰVs��3��(�{&pC�S
��_=���?U4�Ԩ֏'��I�TX����Kv���I��rP�Zrh/�E!o���ȿ��7��0�o��Jɢ`�dӪ섃U>�&G�[e倽����h�1���\��оg-��rwk�P}�Y�lr���n��p��4�1���1��w�B��Բ|jW�<�)�=O6�u3}�'#��C=�s@ƭ�rD��3C�g�+Ϯ}�e�S7m`G4=��g��w]��Z��ȫ
ofM�Ae�S-hk��� C����D��D��F�D�W�=��^af�.�ՀGK�N��Lm��Oh%�J���e��HDe �h6}۶)���p�f|����Q�q+��&$ �M�r�5�� �a��@�,�I?^Z��"������9_��3���O:3�X27���D�l���z4u�r��;Q�Ҋuj0�s�����9�k����6�����(m�M#4C*���)�w�b����c	5�W�Y�@[�X����;Mr��.`��i�*����D�̷Y0�B:`�|v�����ɨ\w&��Ő�`�BM]���Ԃ���*��s#�9"i^hwl�d�����dFC\�:�l���q��]��)�f���ھ��I�����*,T`+�)��/�Z�h�m���[`y�L��d��;z�/��d�$r��`%r�Y��������S��W7���p'���/�fA�����}IB������H
�.���}!}69��J^DϪD�{����ГM���=�����,t���}�jD%�r��#W���+LR�n-��Y��;_�~�, h�q�*݅�W��g����^Zq����kPLֵ�$is�BBaN�g��J���+�يw���Rh�����k�ƽ�!��y�����.��:�������$�D�/	nEt�m��䆌t5��j7�� {p?w���_,o�K͈/�Щ<����{$��6��ft�،&�Q�+��a�M5����*���R1�|�O��bğC�0�`E��*�}/��Y���i�VJ�n���O��:���X��3�.��6b���o�?&I��ExJ�p��Jz�-4i�oWN�a��*��k�qUX���<dycI/i�����V<�e�#c�`���~��mAUӺ�rp�%��nV[�������)��z(U+�a���H�|��z�C?̺dMx�dU�$���t����k`D�ĕ?<�:�	�w����@�D�+՟�i��l�%�b��՜�}����TW?`?pi��d�}TK�
�����{�Ў#vfL�>��u}fcP/ky%��Ly�,��c@~o�$��IZ�@h�[���p�����_a���y���;^��u�Kq��m�Qr�M�v{��jO)�/4���j`����sxw�dj�@j�4���~���*�A|�Ӧ�QZ��P|�j��aL�h�;V5��"�H��D&��J�l�ױ$޺���<�.�̘}��_ɕ�yO��0���h�e�$wZ���o�2�d�x�w`����0H�<��Hy�η�ͨIhr�dx�\�)�,qj��a�y�~A,�H�}���Js)�פT�Bjۥs����ǦN�3^�(���G�G�m�3��ϓ�=�5�Lj#����5V!��u�]��F� �jp��J�Pi�f�gl�g�ɬ٣�\�!Od�$���9��x�O���$$_?�@9�NRlI�3~Թ#�"a6�H�a�/yl�A`��io:+W7�����"�"�Ia�s��4&��黱���\9�ж||&o�패UDQN׾��뒏�\؈���dU����L�!��}�$�.������m�����v�%~�Ɏ�K���0gy�P%���N`�U��
��U�N�k�SnX��N^��*�r��B�ޓ?&TP���?�^9XgVA[X�x�m:
Ȁj$��q�DS�x&�r��+�� �����v��2Y��uC��2��z�+$��6���2<Ό�.�!SW�i%�p�1���^�s�U��������̃G܆���p�5�c��i�	Έ��+�]ذ���:������<˃����ST%�H�)��
�j l�J�ZnM��֜DDMF�;�Ne/v�����9����&T���gJ�w��O$��v�:� ǡ�ڞ%�`:s���h�'3����]��EC��є�a���4�}^PK-z�-����!]DR��e�vI��n;�$���i�jw�>�i|��t떗�x��+��L�YԤ���<(����Qn��gq2���uw~��C����zh6��<!��§�@���X�����S����-�G�%�v@�{%�2X�֝ ��@������{��ʉ[��|�jO�������8e�j��ȉdP�Q<�oRm�u����aT�F�<+��zz�a�Ng�h�p)�E�xL��W�$Vَ��*�
��pw��9^�`8�w��K�AF�Y'�ZJ2�N���Oc�3�珣=/j{�iCd(�����D�FT�Kz6�Pv�S�SCߜJ�����L��f�����E�5�7�I�TF�_z��8���|��R0�E��Z;��WAr=�}r���W��gr�ed<��J�,5}�h���]��F"Z�"���G>��o>�&�d:6�7)z��$]�O���3ϵ�F�Q���ԭ��Vwv�r��`!�W/55�5/lH]#8KWyv�C�H�J=�4� �_��z㛴_֩f�8S^�,��봺X��6 "�k9����i�����(�;n�JB����\E�KB�Y���Gfs����g��4.W�s)���U��]���7O��`@��n;97�伪
��la��aȖ<�\�.~՞�Y�m�@%Q�����2�
F�{�\���2��D!}r[k�0��` \,�.r�_�Q����=�Ԣ�q����C�,��@�YN�!Պ��c���&%S*3�Ĳ?gC�2��I��`�,�!�0�)iX'�le�L�R;�]s��)���� �t&�ZVtb��|*{��e.����{��]�HT��x������4@X5"�^��O�S'̦�f�h�^�K����*�g�/�~�~�3������j��]�r�S_ꝷT��T]�	\[$�}�ɍ	�Fވ���K ���řB�}�˖d��?�w���jU�͚4�yl���إ)����]�r=��E��5�n�J�I�Hu^B��|�ra�K��-�%��[۬?����¦#ƽ�n��
�"׼�lҒ4���9���>]Ȑ[m�I�
�v�!��J��g�ZWOf��r��F����gQ���B ����U�+I�Fy�B���9�`NX��,M�j��o��pgT��C��_Z>����zjˣ��D�.��nZ�4�Ԥ�a�w"�ݔkuA��Tq�o��7,��mT�F$�Ic�����P�<#��v�����E��S��v�L�����M���}���ᓥ"��W�O۷�|�1b1w�����9��ڜ՝������58\{�4���q��Jh�O@�a�:��Ǡ�N��)h�8Չ>�C�������b@h�t���j{#���r�$��Eԧ�΢V@y®ơ���va&�����3�y�z��7hP�۹*�0]�K��KM�A<�W���ٖHb�v���&+D�EN��4���(s�Yb�QUk^Pf]#��&�15�ieBI����ȁUG�a3!�-�C��l��32?�Q����.S�)ވ=M33z�T�K3��7��DR��[u�a�<YE��xU��v(	��f�<H_�ŊS7@��/;=�7�3$���$�>��I�P!����g!A����mu7`���٦�l{�ڵ�#L��	*E�B8G��"뵾+��0 ��9&'���7c��WT�ɐC�&N�L\A�疊]�C�ֹb?˞c���r/��f��]��Q��$�ygE1X��5�z�Z	�H�%I�64��*�Wg��2{iK��f�->�}�A�b�!H�Bs�1�3SW�P|��<]���!Dp��
�J8Jo�{;زV8Q/����_�?k���ʶ�