XlxV64EB    fa00    2df0�ֶ��H�L������X�a��E�菃�=%�"m{��8"���.�F�Ua+z�x��Z��7�4��#�t%.��n>r?#�/ ���m�J�4b���Q	r��o�"Ǹ+x�`!��b�3-�j_�%�rfڔ1�?	�)�$�p �W�s9�����܊���A�tZ�S�<���F*՗�}�2�G��MO�/�h%��ѿZf�f���4����붲��_�֠X>eǗ�:$���⌛.���	���f6~�ݞ�f��vtD�Q��Ռ8��+ر>HgV̦3	ZW����.$�����+���c;��:�~.���Bnr�2z�u���I����M�7#1WV�쑃�倪?����\����S-�ǻ�]N[����/�YS;���`�g�(`;찥�B�9�8ù<i��CU�i������H�t�?���髂� =�x#�S(��e��\�`�f-U���G
A��e���mg� R�Wd�[U���1ӷ�C��mB��b墵��/�=z�K��#�ȂGk֝ss�3���N�=�{��y�B��L��B.~R��a2���d6�w�@���_�\����[LۃܗD��3�lt� ΝAo��^�g�if+����S��q���ռ�&�Q�h u�C?%w��b�뼒�����b�:�Ο'�HeZ�J��n���KӉ�P����
9=%8��W�K��7�1��p����:���@�Xu��C�d&HKq&˪�g&�I!0ۦ�e����c��D.6�)C�%�,������r��u*UHu�R�Ƣ�6�je�Eu�ҿ�s�R/�B�����5�s��Gb.Y�q�}IjK�� ��k���mS{)�_}-Y��!BS���Q�d��i��N�����/V��;t�%{��+*W���ǛY���Suׯ*n=��`���M2�@x˻bS�����gezaϻ���0E�4�jK��3pkw���l"d�'K_��N~w�olK�!v����V(/ԫ{�x
IX*ip<��}��5x+߹>��T
<��I#D�%��#�ą#�c�N�G��sˡןb1���Xw��%���td�Ў�
ŧ�V�e���EV����	��`5�T���� ���E�NO�� �5T�뻃��#(�ȫȣ>���}$�E��ȩ_���oSd֩�$��-bտB��9~��(�H����K5K��57)�nGy4����B��%H/<Z�$5m�B5!{��,�j�͹�XfR�-�Z��~ԈVgl �+=�A.�"R�%�j�[�j��S�[	i�ߜ�[.B��fώ� �C������~����h���v=z�-�XF'�N�87�^��?��$�
6�D�?�m ۔�na:(A�ȱ���$+�O�+JZb�,hP{0����jM~��c!�I+&���w�8�E+Q���U��q��}�k�x#��ۄʒ�ԫE9�	J����z�?��%98�Y�8`C8����e%D��Q��4�C�G��Eh$Ci��*%���{ݢI�bG��a$����Sj��w�5�}����PR��Xa��` ѿ���e)8�᪍4����3�)�w�dz��2�6Ǻ��8S�W��m��2�V��>���zĹ)w>_Z�Gy�D��7W�nث�p�,!����-y� �1A���<����jp���R�E�ٖ�٣b��/L �E�����$�kp\q.l-�5^��t�JR���ni��7��X%��;�c�EX�y.=L�� ��3��/�������T�G��EE�`h?zC���`L�v�M��BhI����.���t���9���=I�))�e1@ `��D��`�%�a��CA��p�v��duv���y��mR���5IUb�1Ne�U��E\�:XJ]�
Ep���+!}�\�ٯ��`K[�L�5��b��$�ޜ۰6=�{�?b0��S�qL㔼@G�Q���3��a[�8���ˡ�����5�˻3��h�%5ׯ*���s�����l-yߠ+��F�{<&y���8�5XH�h�S�*�e�EH5��߳���1�}�)��ߒ�<� !��촧5�6�f�����L�'��!�O<r���S��.B"Q�׬/��^~���0Q�(��#�&[�����>�o�q�/���"Ru���)�� A�Un �]i��d���֐!C����)&C:���wU����2�*v>p�ʢ�a�ns���~!���Y�_����CO+Ւ`��%�AE�5*��wޜt{����r�D1ߝ"�T<�} W���n�}�a�����l�V06�0iJ׶���7����#~�M�Ï��<2�����[Рu��K5��='����M��`�)⁲�t�z;���)���a�x%�cR��HʘD���1r��ۢ���?��ڞ����a�2d�8��o3Q~�b LF^;Q��T��{u�� o�"����w��G���-����;��zKB�]zK""�6����o� M9R^�P���x������/w3����m�:/�$���cW��4��A�a�*��Z���!j��~]���V��eT]0H��2�{��1J�s[�xH;���6����x�SV���0���8�����5�̲�ޓ).'p�;d�,�m�Az�J5��}
?�����YN�t�7��\�O�m�ma��)>�����Ō`�x�%g�bFGt�ߠ��5#2�m��y�-K)��k��e�[�t�:Λ/�d�W���y��@�I�}`6A����1�S�������'C�C2��ϰ�����) �^��z��;�|X_��1�q͏]Jmp���=C��6y+����`~)sk:�v�~�t������|��ēC�B>Y��P��IT��֖�:��GQ��S��R�� �@x}���?2�����'U���H����+3�H�U'�,6���{�&�O$ڞ:�����i�_���MU���A�M��7f���Z0�t��vR_+�E�s�=�6��_#X �:0�����M/��t(歩��]H�����y�A����5aE��<�
y��F��P��9՝	p)ze+�g����BQ����(U�"�2%BI��3iI�|������y��2�1�MkC�̥�6!w��2�?)~I��o�����,��{�X�i��G\�zG"��0�ޒ��d��2�x�x�_���ۣ@ꄲ7���:�-(��lW"藥p�� ܮh �fy��?f:%K2ۥ����h���a�0:ട|H����������^MP$��yvM��֥�*�� �|=D�n$�U�`��)�~�b� � Q�����n�}{��c�	Ż1V�&;l�$hW���O�>�3e��{@%P%d�@?���nk%���ܮ�1�*�3������a�4+�"�������+[qq�ƚ�z(N����_�B�l�Ш<��%ת�}t�j�T�����4����dSܡ�G?���Q�2-����3�\�����r���>Z�n(�vc���i�1����R�7>їO�o�����[�7��a)��G0~v%хz�!����ݣ���dy�,��[�,�-����S��O�4s�؃
�g$�M=遳5Ll�朖���%=a��mM<!|����C�i!�^B�{'�i��˺<O��Nª9˺�Y����}�6�+u���B���>o��4R� ��9�7�g�yT��v�ˉ�����fr�g��(�Z-�w��O�����<�N�ϙ��P�wK�[U��"�)�ǷE�gE=�QVJ���BS�ܣ����������n�Z����(Æ���_��ڸ�h�F2ڱ���rd3�d�sd8���k$�NH�h��������A��pl�n�Z}�������~L����l�g���_��7���(]��J*ڊ	F�'��W��<q˄b�>�ADX$D��pi�q>�`DtG��RĊԀ���p��&鯵(a�r�,k��������X�9�*8�\]�ksU�_�"����g*����m�
���7�"}�#K�%ð����{�����Ft��	�f�IJe?j�}��.s5.N��S�Yw�O$����׷��؆�Jan6�� ����Ta�ō���ɉ�{�P������	��,�8�\HE	X#M�YL����:AlI6ޯpo�l��*ѩ���Υ�e��r�b�#�*���߾��a=�=�ZZu^���5�w��}J�:QEx����?��𠾄/���JL)Y���T�sR�<C�����s������	It�4(%oU�9T��\3��m�4P�$#��"Ͳ�k���r����! �')��k˥��t%X���+
bkC��Æe�#euK�}���a�s����D�c���X�R�b4��hDxu��%�| �-�@�4%��!L�`|_V�q��D�@��4��xj{^ޤ�fO���T�p�Fz�<~���@xja�V������y��4��V_���$m����]�����K��TN��o
:��-r�	��H:�~O(��͏}@�i�
���ŀ��{ r��`��L���$ђ��]X��Œv�"���!��C���M�8�b�,,V�*JM��Q�Z�@>ǃF�!��f�Z^*hݣ�35�R�U�dk����q`/&��m�4>�:o%�f��O4r�a���K帵�B�"��f#�r��� ��%Xi��\ �:�o��rH����7�E�n����?c`��=�n������i_ƒ�a0�ͳ�Ee~!8T�����YuK��n�j]�6>�"���l	2Z��Ş���ip>CB��6X��P�x2�D{'���{����b I͢u)�	����1�<�45�y���T?�`F+�F[�����S3��#J�����6��n�����Lb�Q�{��7͒t�鳘Q(�~5M�v�#�kt�C>�r^���=[��3�4��L�,��Mu��Yf6��t�@��jH'��Ĵ��!>�~�|�qC�KVՔ�h��VXm6�՝��4�8ρ������؏gB�=הՄ��<���:7��`x��z�"ա��r���۾���9�8t�μ��O<ِzvW\�
ѱ����k��rKm}7��lJ�ԋK��&�_�U���U��xA+_=�O��8����ՙ�2�i3���{�J�$��Y�$�R���¢�tS�_y�˞Sܽ pV|�z-�
������BE�q%"³]�A?�,;O9#�����HQtY8AIP�c���������"���Y� m��u���G����h���c�P�;o�4 �I!�(�w�k�)���'kfL�4�Nu�6��'O�����+���SB��c�k��q�"��݋��B�Sh��$�fV�P��|�D�/���[yzqyR������rq��U�`�Ph��=�O���c=��W�jf�B�߹/
h�5!~��uD�9F��ܺ����j&io3획q�i�ށч�yW���L��\U����<*���(��?�@����rIf�:��Q�<�����k��Dľ�ƍU38�t�>���8q���?���.���c�=�x<MS���=���{lV�u4���_nN�j�{gx$_c
�Ǚk�N�]j�8C�N�p9����0���S;�VnC��*��Y�����,�-�Ժ5�`Z��H�>ͨ��m�K�РLJ�6���^bL�2ް�z��������X\�24�,��x<N)�H�U �>�����҉Ҕ?�AJ���������<JM�-#M�.�r2�Y�F͉D�q��@�Ag��z��`��S�"�^����~�5�����D���j��H@�c%�F�JM5��.�)q:��@�M�U�wꤚb/�w�"S�nH���'qJ����d�[-P�_�M_579T�(����&��Fԩ��(�������.g�W/Uk&6��W4r�p]� �7h��?�'G{���a��?}�H[]>�5`�󴗘�.o��V-�*iβ�&ܫ�&X+ߑ#n�;��-ȗ<�%�H�^�(vc/hU�t���2�{ǂK�OR��cskQ�oph�X�}�ƫ��1Y�"1Ь�,ŷ�p�U���*��yR
y���S�o�z����=K|8*���ӽ[L�Ɨ���j�`�k�^���	��Uô����g�M�wa[V��)J5l��yL�</�%kZ�[�l���ʪҪ�+߃tFDi_
��;*O
���%n؝T]Q���UqYI��*��@��Q�.��d�����jicR���Ö	������Ώ�P��)��Dd�01?{�2`�>�wM�ө���7&��p�=A�(����+�8"w�u3��DAL�D�K�w��ss
/ޤ�$��A���ڰkϿ����֥0��s�I�f�4Ƀ�ٵ�=��K40�F��Ӂo�	��"����h�	��)|���8��P���
����TlPi���/%����)=X�_U��W�6�Z�95����ok� ��Qv�Ȝ�u���0`!17���U�{���cr��zBg�n}���vNF�L�´�CF�п~|��ݘ�T��A�+��P�x�	�Nb�q�B^3�u.cU뛧W|^�}��o�S��g�F�5�#�*�`�m���3%�[�{��C�j������=�݌ G����cl��t�(�-�1y�қ��FF��lw���Z��؊k�k�j��eB�,��ұ���4
r����R�b��`(O�<{I�^�7��1CX;3>+Y ��I#��kI蓿�h���'	���[�K�s��Z��$o�ܳ2_��*��}U"jy�r���<�|��Cg�?�W[�d~�&�C\��ƻ����$�{
D)K�8�����'������3�3B���8������O���8�#>Ǭ�S��iaY��7���.V_���]P)s��������*4!���ig�,�+6b��`��s#������iWs�DvX�cf>�������s8G�O������X]�Z������IĔT��6�����r����[��tm[Kj�3PX����[��3�� �z�����Vw�Ȁ6��$���g��>O˫��g�)�`�m���%�����'Y�m�L�����.:��������3��Mk� x�����T�(�-[�c��8�.���ҙ°��U��t�N��cA7��P������ \�#a��ƹ�c���!��e�f�TM_V�s8�Тe����&���-=���rWJ{���.8�9\мzIq���zGzU�x�*a�X��k'�"��э xhCv�a��*0D���/�f���Xt�<.��ًB-�����	K4i<���won�ꉋ� 	��<�����$�Q�'W]�,��W�w_\�	�(>���P����M� Iֵ̎����xn���-��gF�s0��s�_V䋑��3�|�k�@0#бe�U��A{S?�x�jL�@��
D�aN�v�D�ZB�����YF����l�-g�f�.�W�/��nZRB9Q����E�������[���_�Dw
�L.�z�	Н�_uy�l����bt:��V�|����H��h:׸4�fѼ��A���q��5B���g���N�]�?�9L�Dֻ�l*�}Cm�i��N(/V�n����s/�<R�5;�Ay�2�j�����y}7�K���'6)-�+0xJ7�9~v�\*N�*2V��5=�w��MI���,�	V�an��lk0��WIƕ{?���zȖ\V�j�%RʁDT{��UŽ��������րsѼx�%��R���BWE`���6���u�1@�rr)�%��K�Ӭ*���
ֽ���M�������NFG��*��`k5�}Vu�D����{5�[
xej��Wì��� �_AG�Oʣ#�	Dۡ����+f���`�T���ݧ#�C`~Yl��X���L��l��0�6���v��ߋ�����ݧ30����_�Ao�>������-��N�i/R��׿*���箘����>��t�}�D7a�8z�S�^k���:�"��Fo�u,��5��{}�Q#���HK��(X����}��O�ؔC\���V����M�����ׅ'F�v�"8�;#��K�'���@���3�c��
7���;,zP��g:����
j��3J�Ѳ:"x�������]�C��9|׵J�//g�V��7��s�:���$�&���,Ao��'�n?!�x��y�O_8�����=�Zg[A|���%:��k���˕�Qs�S�EZ��p���[)2�9�>���:�&�g`}�
��?�P�=|�e��v�!J�C�c��?��=Ŷ���r2�<�%�L�UYr�=��m��!�uhz�pm���bnj�\�V����z+{�RΖL������lv���F�v����
�ԼTxo&���}���#�Zp��˴����ݘ-	��UC�3�`�(�%�[#.I ���:���)M)��=h�ī[�<�<�J'��-���W�r.�[$X���w������DĨ[�'"aEc��]u\{�'�`�/V�-Lћz�Vj�72e;�U���<�o]��~��n1V����ը�W �K�4<cƸS�ġ��Mnv�Z��)Q=���H�j2r�Wc��i�(��ʾ��&�K7s>gf7�v\�s��^���C�C8��'�/֌.��f#��nw�v*���<�F\s(`��%��7����z�9��ϡ�Ɗ�J,����F�a�1��T���V#Q�k�Y�v1C~�A���֒�淦�ƎW�9�NZ&�����ģP�$��'���[B�n	xŝk�*�D����)T�x���4���Ӊُ��hjYM|��5� ��ʢGtRa�G��eG0�p����|<jT����t��B���a�,�ګP�F�aQr��36�-��|�ĩ���Fj�?k�%`RA�����B���ݗ٤q _s�4pO�_�ؕX��8��,�ʍ����{".�M3Y������ ��߇�}��H�Kzm6̀���U��a��Y��&�p�/����v��<irfL�"
�c�J��I�v��F22��Y��Nt�^9����d��Kf��� b���w@��}O��&�W�T�:`$��I��A<)y$�"�1�'�|F� �	��X�q҃ʋ=gy�[���
����╯ħ������`�C������hn\���i�q�S��=��̚2�:iJ�:9����V�\�;l	vc�ϟk�@&����B*/���u�{IJ��R��9�j�}t.�#q���z���F/���� �z�с�8Iʃ�c �R��k�����j��J�l��UB�&t6�
5Ƒ��D�qO|֕�����|�ϋN1�t��	��x��N��w��G��{�	LB���t@��P��1�i�\���	n�y4�x�ך/��i�����0�{������/�z��c��k���tb	J�x���S#�%���ק�DFus�����MB��af{bq?A������gƉ���-�A1ZwڸP^�>��~/�=�i�uub+S�Ȣ�(L���:�sWr-�d�u{��k�����3/`������3�)�fir�[���4�<}�|�""�ֿ'C�q�����oO�]%��͐Akt��ud�D�|Z���p�8�27��usuB�����GH���x��2�)aw��~��p��[dp�A�k5�l�����ƛ%l	,�_*�.;�ΐ3�#Xq6����q�Оt�`4]䱧�WY�-�=��d�����3���	��#7A4�������
6���&�]Ϋ|d���T�ڳ�In�{�r�˹�ݎ�
�j����p^��[ӑ�z��|
��H* 3�|`5�B�D��5�����ki_�7
S��Nv^c5����Z�� ���^G�,���S��5mK�\�ԉF�|�?ʅ)e�Po��_�p������O9p�K �ɉ��Շv�em�v�����`���F�6���7C�jJ����0f��a?:2<K ��֥!�׾ř�3�5�6J���J����� ����17�eJ*VT��r�[�!EkR^5��`_\!��a�I��羔
Od{�E����/F��i�O�M��6G�7z���I7{!�m^���M��|B����#"1{s3
UĪ�����\5|��Ӫ�۰/�&��n��������8&�BB��������L
Zf}i��D��(t����tV	G���9��tq��})�q�+������nRG�)�+q��6�E����i�$}d�e��Px�3z'��7�!��J3�d�C=N���F�U�B�U�_Uџ���<%%�y�7�J���:�]�Ćc�)�����Q�Me�Jx��$�X��ip��Ph�F-@�v��7�R08�=^�ۊʶ��L��{��RWQL
��cż�*-*8<G��L��bT�^��Mi�/���9o�}��p�R�Z�+9lmw*Ǡ3����w�<�]�NX��9*J/]�˙uF�,f��J{�t/ZFM�.<q��Y%�q֔
�����YGo%]�� ��$u,�Z�w�����~a��R4��u���'�0�-���l�� �v�
Xz���fڛe�$M$A�@KY��I�螆�k�(���򪩽��%�S�{��`�&}�+�~�/:�͎�8DHуb$�Y��l*�;gK�N��``x��30}5��#�`��\U�X-�
Ȅ4T�v4k��9�b�"�Ѥ�_� [�	�d�������}��B��g����2+���AY[s��o��xP�8mDl��_���IM�pe�=2���إ�*�?�u��X[�_(����ߓ�t-��u��$��[�I�部><iު|�v�>��X�jq\��G�?����Ͼ���p�9��V������'�:�Y�="Xˮ�� ��`1�F�9e��Y�"�FZ؎|ɷ_5P�G>��Dǒ�5"|��G}j��\�KW��2i���z�V��!S��N��2��N�:گ����ǻ��呍��c�����D.=���x�F��if:2e��R5�j�+l��	��$�&?�/[�+��V�@$s��d'��6dY��P�;�;�]}�-��J�rN�x��{ �NE���{,�ڭi��b�c哖�X�E��L���M�˫����t�*cy�d^�o���t%��	_�����{�gU�cf��s���m���2Y��>���e��$�`�ghTk�$r�<�Y	,����z���f���T�TA�exd�*���%��i~%�?��=�)�U�'��3��X��;�,�|��)�p��.�Y�ːf~h�3�q�t�6����Y���r��&&����)#�䱞Ee���p��E��/P9U򾹲0R�z1���g�S�I���$��6�֎_.m_��*p�2c��N�����{d�T�(�4���R!8���%0�I"��� <_�]�U���ԙU`(}�p�(iF z�x��l«H��#�oL��B+�,���5��#r+�ky⧕�`Z��7�i5��I�|��ڵ��-6�'�݈�
�|<M��;|k}H�~��]	-�w���b\=5�=#h�C�_ ��m�f�DLf��w���W_�}
��a[�:��Ш��XlxV64EB    b349    1b50w�\�3�i�섴�r(?�h�%|���۫hA&ǻ���q*���E�p�q���f�1�.�Hx�vF��+����&
3��a���.�U(��M�<cm��VY˟`�W�$�`e�����' 2����Q��.��3ߐ
G���[�l/'*t]�N"�1�&��{Ui��x�	c�3�-�M�ڥ���&�W�!�A���\�5�7f�I�f�����˨\Dhۍ�%l�8_���Xŋ����N;D�gaZ�=m���}޴��;}��b��mJx
��%�S�l��Ox6a��1�����e�y���7eo-��#�s�"n�)yS�GS��S�lctQ���D�f�����^�]��>�����ŵ���Mq'����K�1k��DI�ԧ[�Vďa�Rm��*�O��Sߚ�}�<1�{?��gP��7��e�GVT��'��;�kj^���U�#�u�1�}(��$Z��'���l!Y����@�TKL�tHC�7�_P4�I�i��|p�d@��g@���׉i���9�����Q�A�� K������J�t�Cos)>�&��r�.���M��G���Cn�N��9�o)UQ"c�>����S���ܲ��T� ��/��	���qC��?��`h�cj��Z毓��QXL��������=Q'������Ͱ�#RR`|��f�j=�,%,�Yc>P `����wB!*\����i�O!��~B�ɀ��I,�eK�V���
�w���7c�e;���c�/���'�26���֑�E>���>�� �E:���Pe( |�o�h��:���_PSW�yץ�v�6�skt������r�Sp��w}�!߮�>t!��4}�?p���(s�k#*r'����_[�ISEn�&#���T��L�@7ކ=����I�b��'�_Is�+�2�m��'�9������5�5m�i&�+�#+s
�*��6��ƅDJ2v�y%F�ƭ����������-kRH(�%�Dq\��.Y��e�/�U�i�����^Ɛ%1��(��H��^��ۺZ��O��)l�Z��X�cVo]�l"z5Z�G���Q��&x��~Foq�a�"�ps�(��PbU'L�Q���3]g�����z+�agD6i���,vI����!ߨĢ�d�s�f����>�t[(6�>�J�$!kF����&jD��zbh_��;�8{?Dr�Z�Tz�ye�O��~�3�T�y��۶��R��>��{��{�L�˻��]H�y;]��瑶�J�,����a}�: O���f������ӈ�5Q��>���W�D"�Dx�zR�H�>�=b(#nER���H9BV1LU�LI21v���~2Y]-�@<0)
g��Mbg��?����T�����s�b���J{������"��td�o���6��hs��WaS���;2 �ꄯ(�V2���EJ"t����h"=���7W1*m��?#��@�<Ãr��>�sl3�L����`�U���z yms2����������6^>Yin%~C��lD!��=��TGo���ǃ��[�D�L@H�&6w��G�M�H�x[�C��P�����	���`S��`g����T�10d�����J4�e�����]- �4��� �gJ�o�2ġ_z)��C5J�π���j8Q\��h���m&ߛd7��;�@�*�bp?b��9|�ҧ�U����iH�
p��|��Ɩa�N�=���'�{Q�Oj|�~gY>b�?`i�����}�:�|�ջO_O�5�w&C���O
Ć�z��|v~	{�#N�
�`���%q�����Il�r�r$8/���HN���~���o>���Vh�\�(J7a����V��q�U;��"R8���P���/�^-���ޒ�������&y�Vt��R�^��N�y�( ����F" ���"kJ�:�]V�¦I��1��j�F�HKL�T���aX�1m������ވ�e����\�X��G'�K�3�|��I lE�0�\*5����D]C�h�=��M�Z��G�K��)W��+����i�!���ש(ŕ���>u�p���24 c�����
��騑%�~�T�/y΍�Ȝ4z�;���Ԁ�G�bu,�%���i3�ª�
A����iq��1���@2��;����j�Bxb�2�����;�`�r�������rS����u�gqX�9���8��-jE;s�d�Bѥt�c�d���~"�x�
u#���3f���c��5n��-#���ݐ��G(v�-���#��!�@�k#�'X켾W�'���:��<o��8�Ơ<u��ٕ1�����n�TQ5���� �����3yC�xo8�W�D�(p}�&T�g�GtF�C~�YC�R�`T ���6��k�~rkR�d@�cu����j�������A���W��� ��ܸǦ��Dx��G�^W�n�'���a�u�����N��C�b�=�l⥤�L�Փ�x��G���W+�����"Bo��*;�9u�SG��PZ�^�N���b,w��'J�:^�2��r���M=<�޻�j�U���VB�Ji9��7�A���PF�'�Jx=�T6�@f٫�E�x�A��ɁT^x9�Q��j7������S��O���ZPR�4iY�}��y�{<c+�M	�k��D��^�q������y6ϞRm6�<��<�	d#V3)��dF.�Z�͞�y$_;O�/�*�|Pq�N�,�6�?���G'߱�lq�A6��D���djO}A&.·��1p�ey����~eL��y٨�S�wt@1~e��n�W	61�Pb�[��ݺ�m��7�m���J�	-�X�<Ug��z,���*������>�)M���+9�t�b�h��j���m�c�%o�p�jbI*��"�$������ �_+x[�w��,[��vH��h�:�z����z,�Uɜ�@��%+$��#@�Oɏ�,�l�5և�a�'�-V��RU�ݛ�8t�(�+�YN�/��+�U-�nD	����~'PL9I7�=������sԙ��
l�0.�/��� �e�#T��Y��7�cTLa�a�=�Eo�.�W�B�1�X`�dc;�Y��Eۚ�(9��09��98ґ�	:2-b��
c6�l�	Vs�^u�%n�:{k�y��&�z����D�:�Zaa9�e�A�¼ɣ �3t�\
��A������"���Cy�ӿP~��Z�]V��	4O?	��vn��H� ED"�ܽ�)�8�V���?p*���|����N"���a�ޫk\�i_̞_���8�v��t�o�[7�g�`���09Y��nB9���Y�B���Cg��������ץc1��q���E�6>��VU҃�;r�!D�H)"_�3���9!���o͒εט����$OzȚD� 6���W7�mPG<Rnή��酎F�,a	?ñ&EqH�c�T��S�����h}��+;���8��:6R����(D:T�2��m��1
8Y�c�f,�ǯ�X�zF!T6#����v*�Q�A����i�[�}�<��>��R�sƤ���*]ۗ�f��{��K�d㫖�x�|�YXX&c>OF	q9���:8Lj����q~f#nf;S-�@S�4�PUd5�%��DZ����C���B�+�n\G�4 �9�G�	ê�Hʉݍc�MqىtpA�����`"Kt���g�Fԥ�rS��$�AY)�ă��S	uEIo� ��,YA^��[�No�~6�U֠�AJ��Z�~�+��q���Bp��>5����{�حk��jF	Ӳ~�4��'e��>���P�5ץy��t�@�ڶ�N�&�D5/����W����g�>��𚀗f�
�����l�a�t���>Nq&��!ŐL�?�PgJą,��&���P�kh��rǫ��*N��_u���@P�XlY�3���j"�XM��b{���I蛭L�㐌�ݰ�7�K\֒	���m\
e�{lqt!��4�/�[���oƯ�T0~�U�#͵����uc���Ug�trʅ��?j�X�v��z�V=}9�:nݺ�7�'[�	��[QQ�>�`N��j�Kй,�:R�auJg��I�r�'�W�؁��u�)�����0�i����nw���0�y��@� LGմ}��F=-#�y�(��O f#�K1՛�|�iGt�����|f~�n��R�UN�=�*�W�x�g��t!&Smh��3�,�L椆]�!S>��?"�.R�H���7P�-��J�չ��~����D��Q����r��y���ԍ͟s#U��`,�.��T���7ψ��_)iߠ�hD�-h��]~tG�n��T��[1����\	�F2ǃ}���1�KE\a����IOخ���V��Up^��)>,�$;
�I���g��.�V>o�Ţ+f,����ٰ%����9�R�}����G6�U�������ɮ�q4��!$֡xb�)U�Pl�?`k��J/�X��Eh�vK�Sn���;�"'P��'���J���:(~�V93"EWBNN�X*��d���2뛙j�d��i��;���x���$�"Y��qu!d�+�x�kj���Q/De#�Ǡz-b�����t��p|��0C�m��Fr^�Vl�Mg���X�Xz ��;��{��S�Ψ���%�5\:)�N�4ⶅ짦�������Z���Y�%dk����s�T��d�}5�3-xd;�т�B����Mʚ��KI���`��\�ӣX��~�����9�+  )g����uM3t�Cāq�Y�$��):���O����]��>[E�)y�;�:_V�)��`�$�A?��H_�����DC�^�E"��4�$G� .���/����Nِt����b�H@��G�x�y��o���^�ס*��R2�C�k�_�<�G��h�Z��,0V����N�ʅ�?����]|u�����4�E}�먼V����ס�>A�N�E����_Б\r�c��Z���.�������vu�ֿ�	��>+Z�*��-��.E��5�����/v,Bi_����!������^�7h{2���nF�-�
9� ���6|��"}FغT[�^8�� �}��98�(�'��%̝&��sAQl �E�v+,�ܮ��1A��o&W��`A)p&�|J�Ë��=u��h-�d�>z${_�i̘"K��AE�j#a=������(�Zwؗ����%�K�zX\[�$�X|�
M�����8����x`����獄P���lMv������azGS�Ir��̳V��R�r��{�|�-�b��������敁�Y|濎��:��3 b�8�w��J)��H�w�;�8�bj�o���Bw�P�hgz8 �l!K��-�@4�W�-�+O`o���1d�t|�T���<Y��m&�1�x{�5����9V�J}-�_C���]�<���b]���^�t�X>D�,�A��.,�k�D�><!d���E�c�Y�4�������kBH�F�ġ���J�v�1�؀g
y�=��ɻ?��d �E�v��xc��"JN�U�X��<��ŒWq(��S����W;�!�	]��7�hZ q��WA|���}�76)C#+�w�|r������JT��+�]s�bۑ��_�u@*{���Ӹ����-��$�.z�P�yQ��0���)Ţ�Π�fx�N+B˙<b�ga`U������9ja0kJ������x�N�V�����S��溦�WCi��+w�cw�&�~O$O���y�����J�XJ�GӃJbR�����#�}�ЪC�뗵�-��KW1���T�*"j����ɔ[�j�z�^��"�Ш�'�o���<^�t�$�"�0�����'f�G�.���p�##|2a���w�s�ÿ�1��b,�G/bʁ�P�Z��Z�Q��.ok�I}�1�:\Z#s��ދ�Il���g�\2��3@�N	��e�� �cb£YP|B~������5b��_d��c+R�p�7^O��"�?%q�X��K*½���=��� �g��VO�<�R��1��� ��?�x(V����a�?*U����e����hh�X�ob�n\ˏ$[O���/�mW ?%Tb�狶/At���=N�C*2��|��ZZaޛ�%h�3��#�v8e����j(.�J�rJ�ܛ��)��6ԩj1<�Q�I�Z����h�x�$�1<�c[KKA��^�*�?
�iw;�O�@��Ɏ+�c����9���U{���_�E�ds����F3��֠��X���ó�Y���af�?O��O>�k_B���P�G��|�! ���� 01��\zG�XzF������T�o�'�p��6$�D#s>��&f�[�G�t�+��� ��^a�j��(�r{���7d
�r�f5H���Ҩ�&��/	�)x�<�I���=~5 %��+��ٗ�B�6@�b>P�++L�o6�&�K�͋(���ҌEa�@_2KI����5^����6�f"Qm�Fs��Z��#��Eˏ��y�2��Д����H��V�Z`��J�2E�{,T�Y9B�J��ڛ��S\���V�t$�̄kJ�Kx�w\2}'}G����һ�l����<A21��66)� Z� >6��ye.t�z:.5�#�,����%����>�IW��y���܇�#���GJ�q̕28�;QӱTHJa�`:3����a�l�[6>ˠ����`F$>�Z�Wt�_�����4fڈ�"�mwq���M3��,v-p�_��������c~�e�0�./����5�\��`�	^�	�ڑF���?p!�"u6��hXʳ`��;���7���@�`}Z;'D(t��4d:��(<����O�
��������"h)��$0�