XlxV64EB    1b6b     9c0�S�d���Z8�������m�	O�鐛rԪ������Ʒ�2X�o2�]�|,�"���tKv�a[i�I������j�d}�ry�5Ui�В۱vhF�7D� � ��,E���%mȩ��Z=Y���m�#eF�Xt�ʭ�ݿ�}��>k0d�?��qd������@?{Ra���d�#���wc��>7��Pj��;[?�\��M�S��Pt�|���hY�a��J�Iƃ*�D����P���� B ��;|��$xZiѿ�Y��֣�:1Ktt��(@f~�'�-����O}}1z�1��Oz���B	�dH�$[R�WO�2�BWԛ���5f��kB��Ϳ�����o�����I�����j=Kx��ot��?�U�x���1K�P$�U�*��<�{�8���n�vx�lU�������X oQm-�xH+f��/-����֜r4��H��D^}�]��dm�N��Z���fZ3n���	�,�BN��o��T�u?�1�9yWۇ4����:�g]P��i�[@�yF�ƹI;�5p���-�t֢!P�z�������v=��0���i�p�2����ď)�=�}*�~Sj9)�Zc��id��㷯-�ӵ��.wz���t'1�Zq �:$.B'�����@Px0k�>hY��0��v���8ZQRI�s٪�9����R��(�9n#������S�HR��d���87�ʩ���q�J��#bkG��]���ȫ�>`��A()�p�@W�䉣I�(XZ�G����2�e=��flNC	'����έ�K�f��cdf� ��H������{�(�]���8O<�3N��k�QQe�2������A�����'oM �(��s
���e�#O�c���Q��)K���J"/#�\l�� {��R�ҹ��d��C�R�������g�$�^#�*.����n��6I����<��9��
��|���n�J0Ht��N����ޑ�Y�aNo���Pj��ϴ��I=f���v��k 4��F�����Δ��#v53���m����_��� �O� �v�3F�ϊ����-��[���&3	�d�&��V��L��F��p2�c� +�E����s�q�-`3�,7����/����T��b3\X\zg$��݇�@���>���7k��4P������b��S��7o�����_��vJ���D�C�ݛ�@3��8�m��6p\(���K�v�U��JѭQ0�V�8KO*"5����	6�H�a|�����*���&ナE��%�y;�1o��{)�kU?�����љ&qj��"�j����ND�L)���N�2���y�� ��0��G����k�q�!��A����x�Q��g(j�ٙZLOT퐬�:-A���83��'6��sh`����<<T����O�6b�q!$���Q�a��jE-(��ʘ��8T�3����Q#�Ru���S�[E�q����b��2N��o�����/3aX�*���B��1��&Uz���7S�����!���������T�M��ښ�r��%`MK�uw�2 ��>NU\�R��wF߶��+��RMܖW��4��5�;������_�3���<@qq�z_ZK�mqd����D��'
�n=���&b��z{N��!�B-f��<`�_̷�t�;&lI��� ������C2�	Ա�h����'V�`�\qB������6�Qf�h�8��u?� �;�]:�*L�&l#���������Y7�*�'PF��i�B��a���46S����J��<�N�ۻ�z������XW#������t�I��
��u3�� 
�'GM䎫9��~XD��;�[��9�ǜz��@��kN�ç�PR}J� ���4�G���V��45�}�󟌇����Q�����m#Sx6�������{�����g�����g�/?d�\I}'�wE�h_W��2��Hz�CP������>3Z�Pj�t��Ei	��i ��s�uI5l��N<�N{��*֥�u���%c�rN�/^�)���tX�H��l����V�yPw�ߘ:�����/��V�|?m$���p�߽�@񯍔�@=4j�A�9u�Iٛ�X5I.745��ZG�<Ef2����a2����l�`��̓%��vqS�+M��}� �>��%����M�\�ҸCg����?"���%�A�9}�_��N��O��z^M��^f����4�:7-��
C>�����3�na�RGI{-�$ޟ3�7�gϮ�OV��Shk�Mf2%�^Pzn|���vV������'�č�f=���F���^��U�a�	w(Z���&'���L��=�X�I����w���]�#F�*n�{wUVB{q�+�۱N��Ex��KE����ǆ�ozm3�E9"��3���hSh�Cڭ��wE�w��\����a�l����ER��X~�����>