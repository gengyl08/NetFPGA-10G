XlxV64EB    f818    2c90��o��\;E;q<�O�6������\pD3T�L_u�q��\�-�Tk�b�B �V�����)	�5����m(���AƑ�$�V}B��Q�q�с9=̲y��D���4>�����T�
:�\v���/&�6�,���2��ߓ��ZF5���V��B�]}��f�Tl"�Sf6jN�=yb��;^�kr��}H�5"�J����T�n�}���~�����t�+�
�~Xp���~�C���)�,d/ �}_��F�s\��R�><��y�n��T���k����֙=��-W�81m�'6ߜgGL�n�m���*D3(R��%<�S�hFu(X�}(���HЃ�Hje�Ӡ�K�U�*�sǞ���]��n���l�o�epI!�83�Kl���r�J����6P��Gc]��)�-身����R@�g��L�$@��stC�M4 (��h��_V�+�DѯzWz"/�cJ�h��Q����!�<ْZ�b�0�)�p��3{ց���a���BFt�������~�����l%��  %�4��5�V~�B����V�L3�` oO���~���w�?r���gK;	`2ב�m�������V򆪫���}cI�~Ǵ`�-�A䆺�s}���>b��t�F4!3��Hn�loa���M���֌a�=i�Ɨ��mǛT�Z4�8�#��x>Xi��?R]T��H���}Dz�R���� ���!�-T6�T�
ιN�1���$�p;��Kk�&3L�X�J������woӍט͍�l�� b:��g�q�{�^4���o�*I���!v�.�A�ayol7$`��{�5�u���=C�Z�3�w4���>��X�>���� ��r�SgńRl��o8�A���VgN�w��u�o�n]V��gGt�u?����2�\`v�3!n����n��:\�oa7���oIǥLe�)�7M/Z��U�o
��t���/������H�S�i\���q�Y��3o�C<шB���'�D�=0�KV�����G���%�3ǯE�1�/ި�ݢ�����&���>�gm�i�3T*��M��#����?D^��L	��� ǩ!��i<�z'K�X�+��)�mv���6n}�*����X����a�����)ϕ�,���jF�j�,�2����5t7r���qcYZ^�>M�6<�T:$M@���=��-� �6>}�ů���Չob�F�ۨ�S�!��)����}�}%+�TL�E�:S��4ݽbn�����+@Ɏ���e�F-�Ռ��]��zY鼞���z��L�Jj0��?�α/@�τ#Gq<�8�_w��+��ZH/��c���|���QSȖcι�;e~T���@���Hk���Hy4Y���N�fw�B����0��H��y�O^��sM�L�:�Kuя9l;�Fk�bo��d7o*��$J^Nw�:�n��
[�tЎ��t Z�4��t���q�o�CЊ��Zx��Wf=��>��?d�4���Q���A[ߓ1�c�Jމ/���x)Pyȧr%�H���­�)0��@�٫���[m3��(��Ra�D��9-+��'�����}_1�L�%q���Qx��``2�+n��c�=��+��=���$��1�(n����S��=ӏg���[+L[&�8�_�����ן�ԳW��RY
���ȁ��c2>�R@џ}���j瑄:�R/�g�q0~��&|���hK���U�Y#t��ղ�<u�,a��l��<4��K�}����	�x��5#8��H�1����y���ȯT�c�����C�(�A���푬'剨�������u��z����{~ߥ����qh��h��+>R��y��C��w�rF�P�����
K�Н^��ݓZ�mXآ&X������j�A,B�v���,�t{��Dk�|�z!�x-	mSFO�-�s~5S&h�&����>�k��8�󕪆�[�*T� �F��_z�f�B��`&��T(��R7�T�c�XĈ-����53����ɯx�l#��q���3d#n�j��2D y0kOF��������/3�Ni2���	wC��Rݵ��]�k��O�`�y�������L�vv+a-#���2ZB|��W������V�4������'.6������ǔ�G�tN:�(���Z(Qz����_a�ۂ�S
��v��:\�ڄHH��`�&�D���1��;�T3q�[�w��m��\n���
LC\v���Gp�\N��d���]d�}�7����ΏM7D�
���?��K����^������+�l��l��A�tl'l�0��F)�AZ��(,��x>�q����a�m��^�\�Rf+s��<\u)`���[G���e����.X���l��?M.|u���^X�'c�ώ|�PrT��o�5��3�TS�+�N�z�˄�&;V?],#"=�	�=P��j,E����i>-�}� !�����<�����"%�o ˒���̛ ���cN݇�˾R�9$��yiV��-c�>��&�\��������Qrl7������iĸY��f�|�,�ZOc��@�k Y_X+�o��U�@+<,�c%�s�.��,A�F�Ub�j��w�H[��0��Sk*q�v�BmNdY��Q�Y��30B~R}틕J�m���=w��)�5���H� hrg��G��qU��,.V8Z Qǲ!���-�����H��]}�v��.��y��N�Z�oۅ#�C��3���q��P
!��uv���i�.��!Yp�n���ic��~)t�[j��,(�O��޼���[Gc�öjuu P.YC��]K�\�����:~^�fb0��5.˟:A	-����;}*L�o���m�o4���t��/v�l�������nE���|,�
*"�p�l���ri��RK�;�bCj���y!�nq�q�5;��:�d�� \�]�$<M�v��g��h%�_z��wt����y��i,!#��O�5�ن���f[F_:i�]gs�9zA'Y���f,[�Y홃hxqs͓tp���3��1O��},�b//�_Yh��b��7#D�a��0���OѾ�_��L�̐7m��ZY��;?k3����t/#�����6���ϝ����f���3TY�����Ҁ�=>n��I�c����������<xzCU+��i-�@���.d�q ��3�E2U�����Y�OG]峲: ?�t�٩e��!��&9�i�`��	��E�y��� 2pA��,l�Y!�h��2h���>@f ����ȯ}ೊ��(�f�v��a����a!Z�.|�2߬O�x��3X��~)�'��!l�W��L��M�X��ҡ'���\�b�`c���	4\���U����+}�Cd�����e[��]��E�N�v��&�t��M��_�øD���_�gY�S�}�	�^21\��7�IA�9������Q����U�QtX4	��5TIecO�U$A7�X`�33U�]7H._�텕�j,���i:1֜Y�2M�7���RR�ց⨣LS�Z֊1~�1�
�$�$�Ƨ~����]D��I~*���VF��9�i:F���~��:����d'W��o���{2e=��@Fʺ̽��C�ak��c������?�C4y���h`��G9�t|
"M��X1N�U����?t@B}�g�vV5}�g��p��K�c��V�T1�D�;hpT��]~��!�J\bG�� Lͭ�3��'Vٌ�y88�@�������gh�����D"�p�TIȏ�����Ņ$l�&Z�OG3���je�,Q��FIK��b�S���t���rȍC�@(Z���g�K!��NH�
�FF�d@7#�ƍش��'"Im���ju5[t*�_�#�Ic|��I�-�x��bd�ȋ���C�J�䓤=���R��Yn�gx5�K�^�5+�F����U��{�pB@�6{�}""��}�m��]�}5�Z�|���U�tM��3�}*Zg׉�3��t�̔kR�b�Ȳ���C����!�����E��S�jG�$�줙�k�zv9�bĲX�A�'��$��.a���}�&���F�_ς���t@>�����KE":HpO�m/�a���[���A�o&�{!h��8~�?�T����Kj7T�6��Slݟ$£5"�QS�p�m���f��8���^ Mյ4(�^��e'��"3���� �!T1eba�
�w�:~�:���3�&^�'��PQJr	��	A+mŸW�ꟍ`�<A[��w��{& ]�9�UzP5ZI��uM�J+?�lf��#"o�x�V-����Gn�w�z�8���J	�FC��J�ւ2aLa�Lsi��_���XO+�{M���`�;V�c�,��3����.B���߲$=�;�]��5���g�n�%���m���N��*�܇��0��`���U�����KA�7�U)T�����MYt:�2�Q����*T�0�4�1�j�H��79��A���PTE.2��%�k� u��^`���(��<�A���^lb�z�f�	���(�7�[��>m�R]FO D��+z���MP�EZ^,�����+�'<4�R%�+B</�?�=ntg|�!飏����כ�
����+����/����Z\��hZ���5���6^ĪI*1�E�gp���,�̍�r��D�q^�� u88$w�{��/�����B�it}%�V��!�m��Ph��:#W-T�h�v��_��������X-Y� �N����0┒n���{��I?����n�?CP�}�風�c`Jۓ�VwyQ����}��Wԧ�`�Q2�3D�|\sn5�~n�,u�\v~��E���!.������A�Qr��sǦ�2<8�҉`&/�+�.���!�^c/k��t�oO�f7���A��AtD�BB�k�~<���4��@!{�h]��w�H�H�p�0�U{��=�]%�����?�w)��F �0~��P��f�������G����c�����vs��7��u�K�@��s]�Z��-W�Ķ����ֺű8�hI�z���ǈ8��1#@�~�����:�z�[T:4Kvy@��b�TR�|���)e`g�S�G!�qR�ժ&�t�����\F	c�����mY#�"٣�ʄT?R�]ċ� D>]�&���	��l�f.�V�)h���@3ofu�%��H��2���xl�)*�
� o(�>,��?h5��t��픣�˹ދ8���&�t{��%o�����h=�������*�N�N�'�|�x���>������@g���S�I��Z��� �p)�D��UE�Ѱ�������d����;:�d�>�Y� ��9àL(���u����hT:�T(q}a����`��zp�~ZPm�n!ŷ��}�B=�6�/�Ld�p��K���dͯ�O���`F�R@@�DU��|�X{rЪ;��=�m�2�"�j��M��x�u*�>#k]�E�uR�dx��� *�_�hG/JkIĆ�	b��� �X7�n����Iش���s�U-�dx!0L�|g�G E@)�Њv��+w2�Ճ���2��+��Ϊ��a����Hȩ|�eB�q���K}�3�Вyl�<��d=�b�'��!ͷ�0��	�F�f˞"PWdJiڔ�7(�����t+C߃0�K^9�ܧ_��;��ՁÁ5�!QFF�����G�t��$��&_%�CWrϼ"9f�9� Ɲ@��;]�/�Q��6n�'S��J���xȈ\,�:q1eI�dlq}/~�h���Ɨa�2�ZX�FH�c�D��/�W�<(��C=*�f�)�M�å����kA��P�O�g!z�5��%���)����!MB�x��sw�C�fo0���4��2wx�qp�Xh�@|݃i����j%h�ǎ�R\�ٙ�����n�Z��0i���:�H��t��%|Bt4���.��*�yQƋYN��7�9��ǯ�\�,�N}-��!�x_��o��~�t5<�c��<�.�_�<#5�0�׉!lc��,C��c������Aa$�`��n"���������׌�~�m���8�9#@w��L���x��RU�$��qp�5w��`/-�Z�^`>��Ottl�*a8�'�D�Aew�?�XzA:0kD���x��W��k�x�MV՗�˓�ۮr�į�`kv��%!�2J�f_�ؾ�J�,�L�����t�L�^���o�∖�A����?�?�`܇���Ѽ;�'�U���{��D����D�{���d���?��W/s*�|�*��	j�:D�="�;e��\�!!m�w��\�'l(�m��EuE9ˤ?�y���$цg�^��҇�=�iJ4�<��9,m�?��n��|��D�`�C��#���>5����>wA��~ޭ �AUm�u��3���l�M�N3rR[���r�y��o�,"�i�9/Ͽ���f�I�$��"�꾄��8�� g�ԇ]��d��	�~�X)I/��H�d^~3֍c�w$�T���q%<xb�<6�kf {<�+5c0ag��W"YR�a9�5�� ���Z�CՏ)K�׵��g��SuʻO�ߛa��4kv����V:���j��u�~P�Wl�CG6)Pqq�h��4C��0��������K����(a����lq,^��5�¤�tGl8U{Y��c]&Fg�&�w	��"b�`_�����X�T9M��.W���y�{	�g
���'��ŭ��y*Q�QW����Q��#�u�H�����Cl�Ћ�k.�0=�M�� ���eD����K�|Z��R�y��Eۇ�]�q<���t�L]�NOM�<ƋQi7��	��͛=�6�G�3���b��g����}�Ƙ�3J!(a�{�/@��3#�����:�e@�A0"�Z�b!=}q�v�JB���sR8��(;x?���u7��h�Z��8=����Eؓ���r��a�m���V.x��"Ho�(�*97�ȴ85uP4�d]:���F��0�Ҝ�P.]JAp�+3�q��>� SK�1z�!E�9&��ల6��O����>��"Q�X�X�������6�ʁ0�`.�ѐ�}�v�N2��F?[�4�(���Ѧ\�g�l����.D�C�)�yw���w�\P��gF��MbsNJ6�z�ٍ�9��g�����A����������
qyk_ڿ���X@ĝ�� �Bg���iMXB>��U.��������jП�yğB�@ں�&S ;���KT܁�e��5�Jµ͕\�gI
�SQ�>'�I�c�����C�L�O���چ�_��AXJz+�5�bA�?}�≎�Q�cw�c�뫜�c�{lG�ƍYR�ٖ��	b��I
�b��rJ_=�{CE�B���3����p*�AV��8�7�0�e���'��� @�9�J^9*��P��m^@��(ͷa�f��	���Yyt69$��w�+S!������Ûq\�~��)���Cb��t=DR9����>�g��`�BwR����{)�bg�a(<�tW�^xmF`p��to�W���p/�D���R���J"�?�6�9��5�P��+�QA���L���o�K ���<K��Y+V�!el�$�,��EJ�.�Qu��|��j�AcU�{�MiQ_K��[�#_�:C*�(_���_F_���Q�۾���;c5�8��ۘ���O�Ҝ�{{���Y��;�\Xw�N�.���Ǐl�sU����;�#E���8��3&����s��'�1*�B�t�Й��)��*�����.u��Y=ʹBY�r:W��;yx���[�F�ϒKd�&��&oDN���H3�_$$Y��� �tw�?����kX�->ב�N�*���Z"�O��򋸥`����.���"
\��2,k�&~qL������&��b�(�C�)�����Vsy�΋	o���j��uǸ��H��i(�`
��xOz�,0����2��s]���R��V<wU�>8���5���9`)�qV������n�fNwO� �L=�(K�I�������lJ�׾A�>�FA�ٱe�RnR�_�&tw�`�[y�1��x5�l���꣥2�]�$�>�`!��&���z�`Ӥʹx0(2�vt��|dOX���ʅ]��W!�?�[�x�_K�_�T�zUڀ�Fi��c�0��'*�[I�n���}�I�;�|�[ �v��4n�w�6ǜf1Uq���D��X�J��3���K���}C$u�]��2l�~m����/�-7��n��`�3yl�Y��L4�� ~Á�F�_y�l��N�4�_����iUwÈlh���$��V9��b,�)o�sV�#i�$����c?dץ���}�!/4i�G��[B�KtI˺��T�c&$*���{�j�h��i)4�'��<���m�S���)6� k�0PFs�Ɋ�y�=������A���Q������_x3xf{��!֠�]p�T0��P�J�0��~i���ą��N�?�t����QB������ϓ��ú��j�H���H��k?0ƀ��4ҠȆ�!�U�"�V�|�� ��E�]%!��סqL��L��[��Ч���@�*���dÖ�!���R��7
�w�+x עJ<~�ƻ��x9���h$	K�uD��1Ӕ=�5X����?~����2�����]GO��,zY��S��fЛ�%�V��f?I�a�Bs5���.��A���U#��ٿ��)�P.KT�@Z�>���Q^_�E0�1�ƴ'��AUq���j�һm���jx���.�H�YOڲ)����v��:ѷ+r���h���z���KNJ.� �'1:yR,��"X JtO0v�Y��Q��'oD��d,:\��G�,���
 =�7�6>F w�s�U��Gk�7R����2$L�7���c�"���i|n$�d�湊<p熡�cu#(*�sT��xљ��g,뤇�~]0CHm��r��L[E�WKM�P|]a��9:,23>C9�C��`�-關uQ���?]k&H^~}$BY���Ϲ�7. ��R��w�?�f��,t|����~<�IyZI���X�d�Ͻ���&��Z�^V<�ʦn>�~�7��%"[淹`�7�Pu��]���/�萊��G�� �8�쥊��6�>���S.oC*S���h�����5J��s�Ě~f��.	3A��P���T�Ƃd�h�(��˕~�_�&x9|*Td#�1yg�@xd1$ѳ�H[���E�}|؞��B]ެ6p�8))9�;�}F�i�&�ݧ��^Z��$��/��Kb+���ዽ�����c=�;V������I,��r_�ֹ%eySW=����M	���C�㓒���3�����4�to�a�Ah!�@��^��LD�bԖ���*�զ�yvIÆl`v]cY~�$��)J�Rd�.����k�����մ����FDV$�K� Ɩڸ��b�8������pͱ���`s�)y�ɲt���\�[e�87Z����KzM���dweC�&��٤L�fc������,dE�63:e�̤�^NQ���cؕTjdHZ+��@���x������I-��0QHN8Y&=:k"V��ʣVBF�C4�94 ���o
��L�8:\������|�c3������'�{��V&|:����$C<��kB}�Ol_�j$�K	7d��+5߷p>���}�)��E���8�yx�W���#k� � n�C�M�:�j;�H]�]Mt��q,�T�	��~v�}�����F�R�a�o����0��p����U�?wRw#Mx���[��	��f�,4�Q��g"�۩Qإ�Hz?�����N�ƥMTO���8���V�\�8�u����>����)�
��V�5Ƀ��g#�${����Zd𒯚vЙ�����m�j6_2H;ow�ȇ;wddT�.G��zvV��oU���{Q�)�C�����j3kBv���e��+/st���x�q� �ko���($`q�Mb~������󶖸v>܈�I&��7��]IC��f���}�9��U%�;T0�1ș��Z�e�C�`����·f�:�@i�(������G{#[�$-;���!Ƈ�9�,T�ba�����+ڠ� �<��Eo��ʫf�'����ha��W�����#�,���Ť�)����W$�^C����,h��#7N�;+kζ��Ü�ص�R�����������M���P�:e�����`�Y�l~%v�i�� ��^��Fv^BX�-Uu(|;�Q�qN]�6u,;�lN�c<U1(U�>��4ꏏd����r����q���]��A.��O��ٙ�S("�dB�.�m��;�/�a8���c20���aX#P�E
F�;���=�y*/ݮI��3C��M�A8�-�3I�dQ��U��?Ks� 3D�-���!AZ̴�GD�0�BD0ѥq�|;9�(_�����Hrk�sHі���-��`���M��?�5��^"�ԨH�²��A�ju�(�0�K�s���5	l�*s��?4ŭg[0x�y�p��\�w��eq70	��}��B����@���TY���?���c>�R%�ɀ"�=>��F�R��\`�l�],�Z�7�lGn�S�OC����Sg��G>��z?r�A�
�5�k��;v��!�&�ʚ"�3��#H�����]�����L��a�R����D{�7�G�vh�_�{}�7�f�����b���)mB�� d�����{������i,Z(^�AU�ݭ��	�P6X�-�3��R��ؽ0�exG�.a+��D���L���T�D�" 7�`�0�!Բ~E��M����"b#%	��י.����KK�����&t�����NeBݭ��&�N3��� Z��2�nL���2�3�p۝�l��,oak��#�ο��"ҷP�5��d���n��B� ����� s�0����I��߹�ƫ�����)��n��N��0�;;�Qu�Q�_-̌-OU�=���m�	v�yb�`:���j�w+祱Tyݑ�]j�rl��<��sD��-�oCX��Kz�I#.r��֛?s�����k�g7sJ��,��#��W�~��^1� LY��N\���)N�+Y
�}��N�=^G�-2��(U�&䭆(���5Wˁ�EDIO��k��	�6��P#��#��T�U4��w��[��b�I�oІ�N�|�ߍ���t� -"��czN���T��]�