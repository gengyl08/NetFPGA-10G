XlxV64EB    88d8    1f00saf9����	������7�Gw<3n�t�Ȝ�@L�;u{h���ir!Մz��N!�"ޘ���
NWzor�I��5���m�g.�Wi����.Kщ�2�
�N ��=��ጨ���r2�a}���5��lsC��A"���Y�Ny޼����%���{�~;��%_�JL�%e��YEϻ%=�b/�E���5�<8	f4�Fnx IH_��l�'%W�4��L]ht�
X�z��/K�|�MI�gp��<y0T���
���zςn��|D�JYh���cQ
�10^O�t�G�"��|�\$��=d2�V�")����h3| ��I�[`w��"��Vu7"]�~�)� l�[A�-�U�����`i 1�k�lr�x��F�18N��B��`bb2�BH!㤥�Α!���eA(� �zj���؇��~�[��?DF_3�[�O��6��Mp���*�o(�:r~K�ȭ�cP�����B�fo���ǖ�~~��=U�	�/k�����gM�`n��Uj�ؾ�.&4=�6����D������d���<�u*��*��<��<?�v�z!�u�/���b�y1�h�^�l�;+�F��7%��bS�D1�fLU����g)���K�fw2�z���`�5�U;�&�-C1TڗÙ�T����d[�t�6� ���ߒ���7��!�|�ѫ3�Z�d�gK�D�A��	u�h<���߳~�c��C������^8h,[���u��G�j]�)������u�>=�1�`����Ťm:�Ŝ} ��\��ri���E�&�r�%�����Pe���FK��9va�y�����a{���F|Ǧ���ۏ����m�I�qz\<[J��.�(�����x�n�@�!U{����g��Q��焔�ol�o�?E�"���&�
�����m}�vL14�|
�����^n�����������4d
� ���⯡�2�����]�f�Nh�;��6�TO�u�Bmc��s����_zSJ`
���� Hz/���=�+V��/� ϳ*sD�.Z)< [m
/�2jWF�j�P�y�:��gtW(��J}x��l��]�/�;��>��'q8.�Y1~�ϗ�Ph�J��F�0�b�'@�f8���H&�߂�H#d?�I�����Ѣ	�>14o-D���cd����?c��6(��Ō���2�)x�@��VNy�<�/>u��-���p�ͪǈS�X�(��m��}�J����^i���B��F���6��C�fMEd��iݤ�C;}�12�3�1s���r�����8���kd;w)m"��vT�M+��"V'%���[�@C	K����:ֵ��+KY�	?����bk,��_3�~�;�h��&�IA��ב�k-�x������[)�&� Ǝ\)1�sĞ���2S����l�
4<�q-K]��w]��$,F=WՀ�uy�k�L2�h�Q[�(C���;�~j��&u�5��Y���M�@�H�Nc��u	��\��Z�m���d9uK<�7S^D{�|)�\�_��ŦI����i�U��V�&vw��M�W6��I�`�S�-��՞�4���d�����K�6��l@�hQ�,��Hs�s��a�������u�8n���6�~ʼgN��b!#���}��
Q��Z�*�����C'�D�5�Y5�2.����ᨦ�d��R�o����U�li8�%��&�uFS|�_�'/��ƵO�^�扵�,v��Ϗ$��*�D�V//��Uх�˕�+��T�ߊ�"��/E�R�b����@�ڈV3b�u�k�$��=>-)C���@U�Qb�Щ�|���A��f��N��S�r��3���I�s*�Z}��'�y�a�M�,
TG��<��/F#����}���a�,"��H����C_�S�xB W������x����U��E��u�j/�6���6�8M������<��|8X8S0��|�+w��� �n["�a:��u���`���mw�������:�THČ�����Bj�S��V����S�CS�� ~YV�\;3�T�d7E�l\�����;]�[����|��A���F)t�/Ơ�}�|����A��f8u��_���)H��#-�̹���}���v@WEl����=A���`��6���H�W

r`�>�:��n ���,A�:W[�e?��41�G�J�-����>��yĽN�8^�{=;�ۋ���^�l�B�a��1�5�է���
p�����^�-����8�ﬕd�hU1�s"%�/����8���<�h���)�zV�0�n@dW��v4�Xu{�(Џ�R�@\�6�yٺ�|c)�ZBãW���U�Qv=H�7���^�D�O�^���yuͣ]��M�ZJ����r��Kp�f��b>��2��Z&q����#����Y�� w/!����D��s�����c��P���OBB&��M�g�t�.x|]M���>�شU�kΗhQ" �:]�;����CPNc0�3��Q���癁679��4x��MS�ԭ���m�C<d1�w�m���J#��[6���m�^ê�ލCliF���9�o�|��a
��`�r��9�(Μ�u�Q��M�����% �c#�b$+��نhK�,�<iy�ɣf!e0� �sL_|�:���|�����8���F�5�����"��酃KZ��`/R�Ð��Q��i�� ����.�l��f�m:A��!�%���+��J�ͨ_�e��!x���a��k�������C�.�:���5M��Q�p��!���3g4����v_C��Y[��x�=�B1p�9�YPD��oH�M��ߋ%�5E��"F��U�V�$�����Q��KO������ Hg:���r�

�sO��s:�u�'���	�kc)I'�u{'a�e��`��̰��Zva���S��V ��9+��T1�!�����W�X�wś�b
�v�>鐩+IVZ��a�/T�?5����7���<;">&�D�vDI�$E|�&��1
anPD��vH P�+º�H5��Eq^u}�ڶp��A#C�����J	�.�6�%��p�~�gB& �l�g6��3w��x���1��˪l22迩�Z2n�7�I�{��ѡ�)�*�{fw+yHև�J��P1��$JU U�ry�r�
"4�Ԫ��*բ*�	(�|'��
#�m/�^r��Lz2O 7=>�~��;qb��։H���V��-���o�����ѽh~��B�[��î� �l�uq�ѫ�C�z���]���;�܀��^��=�|�~�]�<˅ڲp`?@�6��ޖ�֢���6t��y��z�iߝ�8�O��;���|���rI����8��Јo����Qd��awOgɺ�Ň��˸�^�|��~�lk-��-ү�&; �H�\�-��p��.e��O�$�9i���j?��3��ȕ�K�H�JV^���)�sB�͸�Efj��{�������Ǐ�Λ�*�Xi	�3���<�Ot����\�*��!������~?����3���Ko�J`I����=n�U4}T;̋�I����4�	i+�+zAg�q��g�
�:�z�@�]��bG}�⵴cԹ��*t���9��Zɰ_�8�H㗸��1D��?����QJ��p���2Ũ���Vm��n-;��&��i=�m��!"k��,��D8f)Efo��ۂ	k��E���|��i#ZW]hU����(��S�֖.'Ǚ{*�o\:U�O����">_��*+��Mw���]���"�0_���-�٪���np�3w���r������2iqP7�@wHF�~u/��>y���E.lK��@ÿ&�&&�&_򍃨,f��������G�\)����C;-j9���]i~iE�k$���u5�Y*Y@u!��Ν:�(1z������(�/��vXQT�d���D���lZ��e�pU|�����i
G�s�T�>�%}��`+s�:�fЂ^p:rN�%�/H�*����	DS��^�-�SJ�`dյc�`���]IV��ih��:�^�"X��)
���qo���d�xN �H��Q��T�����(�����tW"�SO��+'O��*���ryk�v]�Ǉ���&�y�5���һ�9�a��+�Fç�s�X�P�f�eW�M�~�FPi�c�l4��Ca}>��*�*��f�?�ޔ�P���\,�����z�?BU1���S��Ȼ�|�ڈ�z~�rq줶a��e��A�G1�YI�.��U:�Nc0�}
{�>����8l�6�^�rRBv�Mk1����������
��-��D���%�"q�>�,��jI�H��P7uR"{=!�D�* ѵ�)O��y� ���ʸ�����Fo�p<]��u���I�ۿz�)��wh�sإ��A+~C$Ϛ�2̈qǓqh��"��Z���yyvC��� cϮ���k�pe ��� ��<���\��<�l�\M�#��n<=�^�ؓD;r�9lCB�0']��.��6J��6&� 	@�[�s�p6�6�'ƏVU�Zܴ��:�+u����Es��pʤm��ܓ�c:�S�]�����Q%���5D�A5��7�H'GY��ԩ [#�)�x��:+t����Ձ��ѳY�/{5�j��G�z�}�2;��;8**�0xx6sE?g�%ߥsOW;��ׯ;�A쇱=K�>�K�,yt��lh�"�uD�'�yCf80N��Wf). @�<S�ݢ\��?m7��ER��~�Yu4��<E޿� #I�����'AK#�u�d��D�KvH�]�ޮ����2��F!�D��L��͆Dq���u�f$��,{{c�Y��x�<���d���*��1��sd�r��H�m����Jc̣�b�R\��:�;�#ǸVn(���f���Ɗ��"~S�`�zAP�	�x�����{/��Cn�m�ոy���C�|3nՠ�f_@��
Q�7����|������w��� V\>f^�I���Df�zε �򐴿vȼ#�"b�Rio8F(�/�r����2"%!*�Ę��@%���&�|�����`c"�"�G���Az�;pp�6�!��bM
[��`�.��L�*k��NBa8֣;g�°��r%j�:������ě�mQ�j��fk��+`0"�ON��L�S{M����-ӕ�D���E�b,����.�$(d�4��(ɀu5t}��C<,v�'$N^��9�,�?7
@$݆�L��^}�����jJC�'3��-��K��ZXc���i��xZ�NG�;YT�h���ͧ�4-uDF���w)�'rk})]�j���>k�ǂ5	`��کe�}���U��`�B	�o�<l+����aF��ꠂ$8�H��Q�_�JOV��Y^��ɸ]I�-�P���a=S�UlUqޖ��6\�/_.��u��YѺ?4��rZ�l��i������'q�;	 �.L�C�<�M"�[zh��rv�g���k�^a��,̸�Ty��[�:�]�mt=��?���˨�}��,�lA8jw:����\�6�������J@I�&" 2�h�����c�#A���բ[5��0��Dϣp��8M�F�$-) z���<�%ܨ^
�Y&���<-!_'��6�U'�o�L(�����)\�F�ODx�&m�W�QS&S���C�STH��Ϋ	��a��3Y����+���)惵h-عf/U(>�p�^�	ӻ��s���go���)m����_]�9��p����~+&�3m��Ӻ��Nv^k�����)b�&�7���'_�x�>�􈖡�w��P��������Cy���yk�p��W��P�L�����zo������x����~�M=D�����mEOۏM�8vZj������R;ר;�b�d�g��ڀ�����*�X)F~�!�֏O�s�TW�ջ��Q�!�.��LV��R�tM%�g<$t��BR�]0�8�_5�6KM}!9~?��~i�-�^�/a[N��H��.��"dQf��JZ�M��د��uL��?��c�WI�����%H����{��d`/f��U$��vr������h�>?2��K�l#CBO�.`1���	�Ǯ�j<i���S>&ӴM}GM�Ű͇%���if� *3���^���O�-?S��>[�^��G��i�s��3��c����W�@�Y��"�sk E�A�2=?K�$�Q�;���n�M����ܽ6���54p|��C�]�v��t�l�o�#��ע�b��<e�:��':ɫq0�m)��Xv�X���S������4+� 	:��$�IC`Qy�4�T �<� ��h�L����LnK_������}P�Ǒ��A|M9�d�|?�^f�j�Ӌ�)��X0�'�D��8��$]�@���xb�l��E�i��<W��`��Nh�/�b$�c�欈��ϺaA���=8�t�|�|�>��pS�瘌�V�v�;��(�
/[��o��ʪ�/�B��ʢ�����|4�Vx�����E#!1�ڃ����ܞ�X��4h�Sie܀y�L\�A2ez;:)�����B�**⎗��#9T���E�K�;�lTI(��z��m��BX�
�9A7l/&����!�u�m3������pc�%R?1,HB��Yɖk7uΐ�)}�ϕMO�JL�p�6���jr�/{������
�A:�_R^� I|�D��)(`�;��RÏ�>"��͠.�*|��Z}AqV�>�\�9SEC�5�P�7����y�L�jV�K�ox!*����N�� ��u����!8�	W��t���}{���Wlv����[b^s���ħ�uv�gra��tE�
�z���s���C0C��>%	4��Vt�z���/�<f3�4�F٬OU�������V$ "u�r��{�q2���+-4�!�9+V�)E?/hQ�Q�:�c����!����#
��ߖ���8x��'g��y-�F ��%�k����/�����mvN��2��q��,�^Fw����w�T�},<1�	9^+`#X�"�v���W2f��r���w����#�!����7�"�6����yƷ��霺�����Nz�c��je���|qo6_'韌W���#40��̗����fG�S˩�S���v��"5O�܇d��{�!�^X^�:��,6K"��`�����9�<;O	U��4��4M&�k�.�ف�O=��mw[m�C%����p�d#|������O!�լ}�l����]��=@_e?��7�S�*�0#?���U��7�~?6-�k��ޒL�/��&�8��?��>@���1aL�<*��(�;ݚv�gQ��gµ�2�uC��k��x.B�my����`v ���c�)ğM�����,���N%߮�<�R���$`-jd��8�ݥ�O�3�^ߐ�
8i(�k+!"3����`��p��!�)�:%\Ϗ �{�βJO�ۻ{>J��w����X���]�S��[yt��4$_(���P�	�+�XQK�H�r��0�OL�tܳ^��7H��1fbƔ"g��䶡ť%��K�]w���=��_�I�(a�~��hksynʶ�$���*��`����Hg��}jnP�59)�(�@:^�E�*Sx��ϼc���!�B�T�?+���ʂ[��W6��٪�]����EX]	<��Gl��<c� �l��������H�i�y�g�,+���" �`޵���S��C7���h�U2�Q�/��������ۼCn�6�%(�Z���7
�~t\�<c�r���B�Z���\����|�!*�Ƹ_J`z�jp�T��g-g�W+rq��E:Zk��E�`*<��=�Ʋ��t�g�t��et?GjÑ���