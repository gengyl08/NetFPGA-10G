XlxV64EB    258f     b30�.U)Qp�iD4pVCu���<�
�c��)K�f��!?�y6�!M6q� rL����l�2H�y�T/�0;+�a��}2�"���FV4ԛ���q�T�3b\����eZT+b<H~F.��@w��hjZ��
�h5�KyH�bA�}����yoEC!l�7�N�)�iB�K�KR�1��N~U#arO��vd��@�0�c����h��Q]�����C9�-]^�����4���<�oK��� ��ٽ^u�o&�`|Y��eu8��!Y,�f�v�
`���QǑ�i�35A����"ӯ|Y2&*
�R����x�9$��9���>; ">�#  ��G��;C_���MY�,�h�T���o��!Bq�XHx.%��uɫC�!�n�Mb�
�$|]%FT; x�Q��.���Y=3vm�93tm{�_GBJ/C��U���`Ѷd����it�]KKF����&���$��L�o�(=F�ˣ��z�G^��$^��
���I�֫�����%>�:T�`~k-��
� 6ܲ�gH����@9[E'	���T�(i�-q,\)0�p�!�K�ph��q"�P��W;��ZW���^���GC�~&Óp�<X�3�:�Ѓ��@��vh�=��JA�;�Y_-�O�M��wS��
xWhjL1�n����*��W�S�`W�����8s��I�G�J/�lz���O����Dŧ ڄk�o��4��M���^��w&��4��臷��3TS���������34��{���D�${���5T'���1��Z�����ɫ��RZ�%�p-4 /��o�pq���
]����Ј�z�1Sd�[���ȡ-Q!��N�e�2����0�f��Mmtm�;���ї�^�UQD� d0�Xp�HN�	\���y��F��?�B�=�j f�^� �&hlo�&n��H`Ta��~r�-|3�؄���'�+'$�[r��/A�$D�%*���[�5�D	,�sI��f̈?���)V!���b�I�}Wt���w��[X���Ie���H����n����?�,��pU)d��r���y8j��g��t�p5�'fȂ��a�aj�ӅH;�`6�#�\��}8�wA��AF�ã(�2%ʻ=�$$�`��+�8u�'7km�g@ ��&�y�L�H��@�rʖ  �3�v���S�?�~��:��;N�7k �g���G�>��Y� �+���L�������3�Y$�d�nC�4ٌ��@�_�CGjLS��x�g)ߘހy�!������l��ŴPyy��K�9��r��J ���Pv�&�(Z`���~u@?id;P%����[�(Om��o�G�,5�B$�i���.t�Z���Xw����B��%c��43���:S���b8z���<[(Ċa`*
���F���1���v�5�mb3#f���f}T�q�\w��������@Q(iQwP}�03kX����)�%���������j�nuNڑ��6��h�@�r¹N��>�gm�X~�����=�nwG�s���΂��Z�C�5K�����7q������$p���Zh3��&HP���-��J.�R`�I��{�?ٲ���U��&��(2����|p��Q�!�����k��c<�:P1Ƈ�v}c��Ҧ�N�Eˀx(���Ծ�яΙ����n�� ��ЇAh���Y��D]���ϳ���� |$�+A�M�+���[�AŚ��|�La�4ܰ���������b��z�6rBQ>$�׏��8Z��Ѧ��G�$��D������Mu�?�xr�Hm;>��Q�-:�e���=�.��vk��%�s=ij��4�A�R��"�a����R��~�������;e�����������衱�S�4e�>je7�w��4��_{v#�ddw�UL�����Q�6��@��9n&jي�7�A�'�AB���Ȯ	��EX��4� S��}w�.�v�¸��}r�;��[�0=Q0_-{�(5SR2[��Kޙ�T	�����q�^t�AƱ����a sm�P	�9��!����85͘�C�Z����@���t-��*��`V�]8/�Ɯ�i6�9G�+twD�K��v ���ce�knݤ>AAx�M��s�ܵ�^`���o���A�\��m�B>�Z��	H�x��+�ĥ�;@8�΀P	���}|����P-"B����U�� _5���9�X뙰kw8K��S�+���қ���@JL{J�hX���Ά���𖧴�%���;���(˪;�)%~�}-p[�����\�O>R�?Xj�����rC;���Yf�����^���y�'wa��s��H��05�����XZ�^�N���(U���&��B*��2�g
��ھ�j�{ۚo��x'P�HW�B;�A)��RU$�?�P�ω!j�c�������j�t��k��d2�1���f?H��1~ʝ�݈���Θ�|�!��(af�`Jm{�n�0m�V���l�W�T�tT��7�2���Ř�S�.O�
y�y1�7O�jP���
>�u�ӆ��@|��d V�R�~ɢo����Y\��yY���{�i��@����K�u�����Fl#�����w��}��\9:�Y�,�����u�=�4j
�-�e�3`���-W�^�~��R�;�J�;6cj��B��M�SΆ�[�`�q!�z���pb�5���ٺ�b6�4z�B�� �1�},��@�QU�)�k�O~��j	�yݕ���-�F�3��;��94� ���u��zf�51�뜸ͣ���>3c����g� �yS˻���׸��H<�e9