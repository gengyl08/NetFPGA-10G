XlxV64EB    1ad0     9e0��7a��a� �`/�0ԝ]&��қ%H���xr!���T�8_��LE���'J��g	�0���(�u$ ���I�k��V�R��h�*�zE�4C)ZL,�{������A�T� ,>����S>,nE���V!���؜Fu�#�v�4ܽ7Y�#y��+q����ul��?��G�2�K��V��QD���j���k�Fo���gn]$��;�s��TS5!��uY���� �UT�-$�0����ܯ�ReF�*Y�9���l/�wC��u���Mf��:Y:!��������ݜr������'�v�#���n@׸y����w�A_P;���vw��{�Q%AmE�<^B���9�m��<�vW��O�f���e�P��fI$��q�ۄxyy,�M�k^ѕ�P���d�t�Ľ5G�BQ"c����K��� .�N|ʷ="C� ��א5�ѩ i�"�]��D:�Ŧ�Q���!�8�FPM:��X^��y
�5%e����O��h]d%=�K5��fOi�90�v?#�E���Pz��L�﮺V�/�&�т��K��Ÿ�z����K����Ya�/�5��z��4=[NKZ�y�%�F!ldAKG�'_�[$������inrDJf�T,�+�7ٚy��.7�S����'!s�.�����eB���4v����}�w/�����a�Sɢ���Ȁ��;[T��!}���l�ɰ35�d��o������h�e���E~X��p��q�v�r\_*0R�P枣�H��������\8�����@Y7OH}��~tl�Ф(��b�t�'��znU|�LM��t{�%ß`{j�w���PJ.������u1c:�^�T��m���fߨ|3�_+/����"1r�/|Y�FZ�2�l���MYE
qLѝA����𒌥zq�}ң��j��AyW����S�Mh��� ��{�*�۔S?4ЫD!�g��N�����͘ �?�Q<w2��L��x�E��]ߪS:�-�r̟`�=�����k���_��`m0�&O����������ғ�O��
ˈT#0�u<��G{&=�S����i�l�*��<��O_.�V�	sb�S,�	q(���N�' *�x=�'Z�Uj|��ZA���rX���E����$�ݘn���W��)��>��2s�����@u�um
F�)�/��"��h��,���i�V��e
�;q���YلX�^*�n�`,���7D�lt悽i�!�. |�	
҃��D���˄��0���ފf&m*�U�ø�N��{by�;r��D��jՔ.f���y�:��D|���a�uP�G���,���.2#�0�ڌ�?�n��oLe��n��0
ے0�'C��
lvZ�����ZR^��>����l�}��8_�"�w8�"���S��.U�,�r��rѳ�������˟B����@Q�����1,�s�!��F�W�l"��q+{j10D�~ss/Ϣ�����b���p��՚���T��oAIM7=O�Ն��(A9��R#���sX�~[��1�F=N�z�[쥢��Ȃ+�5cC �
<I��O7���څ&SG� �V�OmEZ�J�U���� ��*���D��Z�w�l=;�L�������c�lᘄ�6�`�������W���yg
^Ȩ$9��Z�/U)������f�kO=|�8�.���8
ݢJ�vi�J�f��u�E�}`��0��@�>~/�.Y7v��h;? R
��|�� #F�zP��N���_`�/�ϢW�>����� �������z�Ӝ�g�~�f)��p�?Fip�-�7
�?u�Z�A�`w�6Y���j��2���.o�Ff)�{><�n�u���w�Kj�)��h@�M��0�&���c|R����2Է��	H�#9gD���$�uՎP7v[��H�ҙ
	����+��;�]�p�j��r�6V����C����>s��\�~�외C�W"�NzJI�QE�{�Z(m)Jp	��H��	�8d�͕���P,���#��ړ��>��2�";X��7lu%���hyeӿ0��ƽT�ʹC�y�Q'��G�^Wu�)��*�J��2�h�5{D��]V����L���YF��vU�5C�G��n�$��W�%C9�.��uV�p�t�l�Z����� ��N��pk>�b�^���}m�̙=Pb3
�9)\�F�t�1k���G�9RH7��2�l���\u�s�=F�nN���(�?jT��-�;��d��R̍��9<_�%?�/'g�����&y�߄���/Ck��rw	�5��n��n*K�]�m>�X��vD�qn��.z�^`�L�%w�o�a�BMR/�3Aݑ�=���.�9Z��|r�P���V�MI��l;��s)��������	�6z�52aV>D�#����[��w��f��yVv��wH��t��Da�|�z�Xz�yՊ\�K1�>ԎF����}�3�nm�������