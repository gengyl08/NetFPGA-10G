XlxV64EB    181b     980��1����4��=�;��`��ߥ<�&�gw�'F��w�'�h5|��2��U���"
��63.d�nı@aY\��л4�dL �G�n�������ԥ���\����y<�-%Bh?�u���=.B`��m*1��n�RI���-�'!W�Y�^�"��3��W+�#,�7;�i�:ĩ�.7*Xs�C��h����8RE�L\di+i�"�(l����$�Y}M2Ŗ�h�c����WO�R觜y��X�4�N�Қ849�~��o,!Le�,-��WN:��O�jOv�="W��Pg�ۙD��-s: 
@^f4+m_�������d(��z�O2��H�bWW��&�v����N���r���A�N�o���m����'(������;agϱ�
~�>����g0#������"�����%��3�?#mB�Ț���g�l����i���A1��(1�Y���h>�/�'��mc�A���q4oP(��.
=��&����W�= 5����Ѣ�ăX{����y[��U 2�Y��A)-��A��z�U}�g1�]��xjY�L/"�]z���Ʈ���>� ���H���-�a�6�Y8���hα��"��S-s^K8JU����bf�1�]�96y���@𐌐v�!��H���;���	��o��l��K�>�a���3���Dg��jB�Z��s��Lo�@H����4>yr4�kŶ:W���^�b��T�W������"��;S�}��C	�n{T:6=�y�^3P���!_�mW���I�y`0����z\�0m/��1a,E����G@�;go	�U�#����]���vv(��/P��`ߚ�i�:^���2����g�+.��h�lHu��~E*KF�dmC���&3���3���p}�T(�ay�q�NJ�j��,#��2���sia�g���ë!���@�-r���<
�.�l�zU�����͝nN@����X!`ry��]"4����eSi8�>~��̕�>�p�|U��@C��ܙ��ŏ�7��;L_,!�G�1�yI�_;Ŭ�RF����J¼�ӆ/(		��!SC���K�L9�:wa��C��y�%����fh@���%W��z�/W;2d��r�Kb�Z�o�O��gw���)�kg����"lԒ��}��2s��#>QD��mx��1�&n����@uB3u �2������j.V9U"�8�v�&�-i�6n�2G��n����.�mľp�ORZA�9�FT�!r��a���G�&俢2fI�����+U��d>H��p����&�U�cqr�î�� }�55��M��k "+],#}�����G��~W�#)r4Z�<ن�t8ԃ���:��j,S�v�sa5���}e?t�x�&_����%�K��5(��4X�����2Zf�����+s���3�O�,�b�x��yu�'�y������J��v�H�/����ԼR�E����������&�\�2��ܥ\��cN[�*X����?C&�%�x��� ��Z{&W�J>H�Y���)���o��&�YF�tJJ`N��X�f0��b`�{eO�~�9�)�m��(�بj�k��p��[%�t�Ye[ϧ53���C�O�����ϲ\Q�"�F�V-�߆�o凫H0J^߅,�͓-">$������t,f+�>P&�7�z���-��AW��҈�rf���ƅ�Vlms�ꆡ~ X�ϳYor��~��a���w�tBY�d����K*�NB��˗΅L���v�մ�^b�N	�ie���7 �.dk�sl�Ɔɗ5��3c�_���1�o\���:1�*��P����12���q�4�@�$c��I�7`v8-D�E^Ht�%���I-���j�,���<�&��ni����|�^:q�EQ���9>{Ud��iR5�\aZ��s�����ιJM���������(�����r������ZK����$��[�A`��V���sJ�q
�QB�b!��x�v��3%	v��#��G���� طY^���*^���݌�֌��1\UA�#��)QoU�ig�B��[O����=q�J�y�ʤ��ï�P>�7\��LQݎ�ٯ0ɇ�L����hXl�^��>�g�
5
ݯ�V5����`GP�g�8��u��k�.X�^J�cn�v�Mr��b�����o�#B�n�,��CZF�"�[�����sW�L��H�OV�]��le����H(p�ti�D�X�fQnJ`��<Z������f�kdX\ԫ���Va��|�bJ�7×�0V���+m��ys�����_�]�)��r�����	�t*�ΘN��/[��N��^u�]Ҏ�Q:7��3���|����V��d"����