XlxV64EB    17dd     990f|!���v��h������+�+ p�+6C��c�g4�[��|U,H�p3b#q�ea���Ϗ*��Ԉ��zi5����o��n�1��+�XO�iP������Ƙ�DH�1j���5��,��T�tk��5�C�c`�E�j)��"���cc`��G|�t7����Ha�.�7hҏ���3�z�Mi�z�%SF}�j�Tl�O��}��=�d)���ꈿwt�D7�t ��Df���� V�y�k�56J����ܘ`�8�s1`��4(Y[��#��d��H�5}_mP�*��x��$6��n�]B�x�������s³�&���q:��o�F!~f�z~�<����' ~>�#�W�����YŊ7�!������L�k���&;�o�+�-y�p��T%�Þ�����J�D��a3��p��j|�0|��o�[W�y	h�ܚaӘD�?%�C�xp��PŘ�SP/X6��f6T��h���'+��[�c�=��zZÖ}in�;M�&(�9ɜR�fu���i�܉I]#F��'��y����&#@eP'Å@2�v���{�|�WI�˛V+*��r"9�Py�B��n�m[2�8mv�����5��6�Ŀd���$�XyU�i�D6�;����Q��d/_��%�C��?1���	F�<{BD�6�F�qf���Kd�Lg�/&�Q�0���!������(M���C_�~nt�h�"�H��<u�ﮘ�x��p�����2���r18�NW�{��j��b��#��I�8���"h_:L�v�Nm��I@�vE�^�u�\��dG�];;�s�\w��Y}�#�g�U��LXvxfy�guEӝ�wӽ��SJ�\l�_�'h�l[��3�4��Ѫ"�g�}�k��I�^-��{���u�
�l�	=N�B��2�>!c�Hko�S���r]�br�68$��Q2D��(C���aO��iu�ɭ�g�O�X1���l�K##����N^r:JBl��Pe8�`M�@+�=�jݐP�(�{�=��+�����4��PC9}КTt�$��?ADP	��`jN<@�H.z��|YF�-u<#�_������J"}��	�r����h�s�e�}}�Z+���N0j�(�>��㩱����퇢\A�	*J�[���E�?}0�'�"�z��ް���΅��� ��r���Ӕ/z�	?�oo�P��0����g��A�ޅ;�F�i�#i~���N	/~o�w���� �b���'V7�@��U�9U��d!
�V�cR�r:�@�'�:�����(��7Z
T��x����l,ӫ��f�)��&g�O��:�gw�N��hg�鯬�So?���u���ٿ\%gZ!׼*56{�&�����R�)so�&���b/��!8������И2����q�H^�(�]#��72�2ʩ��ȋ����+ۦe�
�r��$z�=�W=�T���|��=H\�B� %�j�n��{t2� u��ȥ<+���v�.�Fr_�ɼ����pˑ������Kf����R�O+LQ�<�1�����5
���3�_4��DR�W������[`5�V��[Q���a��wO���%�4��[��?/}�;%��zR�@p���9ś�¥�=�Wi2ƫ�6U�#+��gr�s�v �ړ2��cJR��}֣�ϯk8{����2�����N�T���]i��>^B�ib�4�V0c�=���%X�u�r����s�� �v�����|�3�����kh(���ٖY�+ 8ȔP��Z�U���HlYUų��:��8�Ns�>��Q�/�F����P6�d�߯aK��ڹU���F��D�@�Twd���:UC7?�(xyc��Һg+�o��kM	�`�&=�������!��2����u�&t��> J��Ion]�����؞.1�}nt���fy��˃�����x�������*c�9� �����Z��&�5lM�:?�B,8�{g�� ���4��^���҃Y�fo�=���w�#�.�����f[W� �~�Ĩ�@r�!Kk!7��9��b\0��8�0`�m��m����>�i���ƥ�I���a��b������+��Z%D��,5���*/\X�t�Fx��Q�y�C}�h8�>�񐢗+`��� P.�Ph�0���>���tTi���Q��*���#��F����D={�i�|S���^O��aa8�Re!��ǖ4T/���O,.�덃@>$�Y�±�����t�'l��r*����8=��J�D�H�b�^x������@k��`F���a�������)fʋh4�n�j¾�r9���܆�$*����N]�t=O�\T�FM�}�"�Ǌ����c��[��V���
�����R�&� ^�����9Q�ۑϝ^����(.�