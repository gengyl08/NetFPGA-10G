XlxV64EB    6288    1710�����&d�.L��qA�c�
'��d@E���%�k쟗�:���%{�B���I����z�U�F;�:�n'bw"�&����&Z��&�Ҧ���A9<�zGh��m�bA�&�BEpX��R��C<��͟)XC�3�kV��#�m��'�@���<�+í~��#��(+q%��zX�:������c��"K�E�r� 치��9��㚴;�X�B��:��f��x�8���νR]9v�1��;X?��+ᖆEa��{�:(�>�Q������钪h�	^^���ZH\����O�G n�[���N�=*}A�Rz�'k���E
QW&M��'(����D�1:?�a��E:��Y���hV� *U�e�H)��D./�CU��@����:�9��t��v�u��/T�h�F�(A�[��q��uN{*�����3O�2�6�T�����(1����3S�3��Ɛ�%B���a�i�c�Z�߼��s0��9=z���3_��лDi����c
��yۄA��g��C���5J�vti"�%�Z~ ���]���?m>FM��&����M�~n�l$��x1�;�T5�W��!n�Ԥ�MDj�T��<�MX��aH1�(��GM.�ɫxfY5F(_e[���隥�N�p�/R���0%���+e�W��V���Z���w���3�N���gS�v�K�/lYO�V�K�ݕ��@�H}k,���������[��6�VmhI=���~�+\�lZ��Gz�-�E�s�p�9������VVss�_���Ƣ��B������Ak�t0a��Ӳ�s-���y�����^&܊�-�p�v�S�����	aŞG�x�k�G����GW���T�u`+��z�%�M�B�G�jju�?�1���ᡟ�)�Yp���|����f�B����ď�߾X�i�|s���+�� �Ґ g^��y�����ZI3�!��%cC {����LQO�����LQq9+��-h�oy�X�M��|���^`���&ߵi:�J%.X���� G)����U�kD�gl8.�O�%�r>6�I|���
L��|h���]�{!���ט���L3"�ԅ��@�є�u�Pm5�:tD3����M���"�㲅�\^Ɯz*y����ɉb�f�Kt���lB��(0Q�B��SF��Ր����Cs�J鏭���co���Ԟ��K�u�]J0��݃�j*}�QId�ت�g����L���R
�9&�w���� � �\L.������_[*���Ms�*����V�ʚ	�8�(5�<̛ҁ���ϼ�OD��U:X�p��1�N��ɬ��)�]Z`l־g�7/����7����c( �����繡����j�k�Y�SC(����)�U�oM�Y����j�-�Ħ�K��@�R��e�q4�^�p^����-p�e�-wU��3�m�t"?_�*�<o�X̏�[2^��	�����b�����6+o;���ꨜdl�AE�����X��+���.|/qE�������X�ѻ_=W�-N���)c���y��=0�A���K���9�����ZZ����v�少T�Q�O�N����W�"՚"G�i&�A��v��Q��ZB_'r�Y�aD�&$U��2r���T��c���!��D;р�G�GGw5���uvAľ땛�}�C`/���i|��  l�%j��s;����l5��t^V�Nx@g��=[x���N>�.f)HW_:�ғ�f*��yU���5MZ4H(�Ȅ��ŝy�<D-���po�lZ(�ݨȩܶ�Js��tKDF�#5��c���_�������&8o-7U����D�i�7��6�W6(F�s|F��b�}�O�B)�~t
{)���1d�D�,}�q@��g�h�2Y�'���@ b)��3���ѧ��#��4�W�{/��c-f	Ł�uxȢ�s)X*���L5.V��K��8_�I���(pr��P�|�%�|��ՙ�]7����!��8I �X�Q��$.���nr�R�,��0D�٣

�����+L���x��?�H���|f���[��W����!��FyD��v�w�tact���WYx�C(ƝTD�2���Zo|Dl�Sd�&��a�w�;d�D+hRá�����X�Ëڏ�L~T�tY=��QH�w�Q����wi!C�A�@��D�j%0�<.��Md�L�f)�Z���"#�Yx�c*x-���Ec����h�4V��n�p`�i���`�S�E�d�v$I4-L���R��mbI��3e3$UABbS�Ͼ�K�=�@5�������*�>�x)y~nE�r��l���0��Ҍ@�,���ja~L/[�����l3T�S�i.�OA�]GD1Q����o�����(��Ī�t��� �l�f�0��T�Zu��5���NJ`j]��I��_�1�޿v�:TV�)� }������#R���?K��L�>˽�b�OICEز�^�3=K���W�P��j$s^f��࢏|���4�&e*o��d����'�4i3��b��p �����<��nz"!�� ,<䯽a�5�JȖ190���~X㩏*�=},� �yo"ܚ�w�5Y�ߦ����5Ɵ�5����?��`*������Sv6�GZ"�g5����U1���1c���=�m�(v<GH9`�.]/��(���5n�Af"a� 	��Eq'�Y��ۄ���|gF�c?4�Y:�����$#�E]�a��f�V^�.`��}KD(�1"��LB��n�������pٛ��j_:��/���ĭ���i��#e�X�k"�����'�e���q܎cβ��c�� ��2�Da�g"S�%�v��sH�3�ȫ��1&�dGޒ���y	�����W7���{�"Nb�ބ\R�Z�m��Oy����|�u�=*��N�����N@K�3� �)�um8JEg��_���C5ZQtqBV�U���%C� O=���C�n��#��D�V(9Vw�v?���e�_'���E�g@��BI�'��8!��p�@�	=�owM ��	��5�"���&�CJ~����f���ݛK�?�bIGg��Ѕ�`�}���w����&�۰_ۂ��)&�H��]�G0�ٕVq/VM�i�s��1[�*@e��^v�0b�H.?�Iw���̂���:s��M,�������c��
VP8U�aZǰ#m��� �M&@#�ƥpw��w���,���s[������$?'daǦ�w��7u͐��!�&�/�4�G-���l�{3����o�<ZM�Y.�ig�sZ���\���� � �䖹������z�:=�X��ޱ��n��z���'����p9R����u��ZSsK��<�L
_�-׾���l�Mx��
+�@��f���q��ߚ~R	�f�;U� ��Xg��� =y��uU����Xm��J�5��2���� �	V7&�^b_�I�����t�2�N����D�Y���  =c�T��HQ�~W�Z��nf&?���{�h?�d���-1���_hIX����\�(�a�c����>��<�3N�]w8D���Vʹf�5���Q%?A;Mk��_���%�Kf��{GR?0�i8���ɥ���|f��2��^�)R�Z+���ӭ�3���<S�<ƇI`wIc[�MHm�f,�ɳ@�sD�m	�?��os����@3��S�ա��9�K����}"6�J�kg�u	��N����iϲ!�R��%��̠o�����R%N^�
}�s���E�t�65q���.������DQ����2DTVĢY}@�\���q��tN�I�tdiN����;�hu����+��:I�̰��ؗ�K��҉-��#q�̹��-u��O������Og�k�G[�V�
�a��D\�I�yX�	#	vŤ'4Ts�O�Q���4˓;��o��mHM]�~� �����6̏]�e�����4�����a\ P �i=J�K���[�����:�%|�l�<'�!���B�LbrH�*L���TE�棓9-f6R0޺�6�)e�m�FK����PzirrU�~���`|���D8�����X�stߴ��K�?Q�-�t�\~��q����Y^��u���go���?�����r��O�Ss8^s��\��h6^KC<�_}�0D���BY��DcZ�mS�����x��p��P|���M�'E��!��5-P6�`��; �²��l��N;�f$V��)��t���+��,�	�u����ߙ历저e9��>� �����..:90�w��<�M��B})u;�l���M��av>Z+Y��*߮ف��;��C� �¸j���i��S�v�g���lpQK�|�y%��ac��d�:�T�̰����Z��u�#�5S���7lˢN^�o(-Tmԣ��՘�ˢ���3��3Ր%�1�|1!�d�:N���n��ĔNĭ8�u�IVݶ��*K=,m=Q�����L*:�S�Оi�5�xe���xn�A�C�^�:�L�����KdEfTb��;����Y�n�մyTr]��3� �o��F��{Rͺ�z6�C�p)M�sU��X�x�ooQSfupf�}��{8��a��I�Gp[��0B/F%n1�\'-n�>��9k��5��"��o	V|̙v1fW�lӻ�eE�c�݌H=�ѕ���H˛���[��w2�{#�w�H��h	C5�!�f�%�L���`�&#)��� ڑ� Q�i\I�\"ƽ�*�Xe9B����X�ިA'�'��%j}����A���1,l?�#QՅɃ�Na�}"
J���Ȩ`���Ϣhd�~J�B���&�(E:�rĚ�M�^�T����CY�F�7���/�M���yg�����I�e�"���;���F����`R#��u��*��)|�b�ܻ���{�h����u6�����!S�eY��?:�v;��wE�?A'��vz�G��xh��L1���B\*�BJ�����*��Gx���fLQ��>���T��Ze0�'���1;��<v�+���n��S��G����a�x��ǌ9�6MRK��Tf��������.�-ex[������?����ǌ�&ӛ�Y&��U��gw��c,��Nq@'X̷q�%��G�c~������@�
��l�P�~�	� Q��8To/ô�R=�,H��ʭ�\�:ab��U��fW=EK���rYE'��E�^<�j7t��cb�{��$��d<u�>^�=����}���1��0W�DͿ:MRe.������/[��!���k���t<7HƳ]`� [Ȣ�4ԁ1N�Z+F���ߟ�;7r{/_�4�<4E�P�֍�~mU#��O�ƽ�+�?;���e�/�}�}4�٦]HI�2덕\Ie-�9�t���]&�LΣ2�)q2��5DQؑ�&���:�H��������C~d�J�� �X8��Rp_�[V_RE9��{��ݣ}��w����۷ְ9Zʬ�@.���)3q͛�"����cbh��ឣh�5�ٵ[ R��ׅګ��+��2���2�6�G��umA7ѵe����)A��{ݝT��9�W����Q�i+���dL��W�����  ��w�fH=ʘ��uV4��Dْ�=o�3��h�#�"Rp�5�I5D��F����* B�f����f{y�,Zӫ�W��ݗ��k�F$���\�������OmDZ2>ŷ�Mט"a� ��Ղ��w�%�����R=�Yf�xW?�熟4���'���a�d~������z��*���nz�I/�yg�������e#�����5��۱h��r��\��j=2�Y�~�N�h�����G+�/+