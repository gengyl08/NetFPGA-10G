XlxV64EB    2b47     c40<ĘJ~�3��=�D������
�n�wb���RB���{iO�����{'�=�|������}s^i���u�^��Tb��苓Z܁����@!�]R��r}�|ܩ��7�F���\�>D4!�"�c�1���0C��%�!���>�gR��ݨ?�@�?�!�Cp띐F�>���I���=Sx��ÃoP�Qw�[$��ֵ�_,�!�/���vՖ����l�4^*�����3�χh��!˽����@�<7���8���ar�e�	�"���kjH}wZv��1+O�ض;{Dc�!ql�W��0�Wr�����e�ӕ�u��M�Y���`�&���mhV�&$��9�4�&��	Lظ��?�%�:��n�PL�A���mN�N�wkȢ0�g��%���7��ޖ���8����~ͮ�%��$b}���`�����e�8�c�*�k��{�Ȩ�7���P�r�!����� h5�R�f�ʒ�JzZ��@�{7. x`wj��>fM�0�)�]�=�����4z���˅U�S��3�b���>�;��S;�>� t�mG���[k��rw:�gx��1ԥ�" S$A?������g>`��S,[�黫�wK�zP�S��@�NOv�5�x���އO�W��w��9�m�W%gU:A-ˎ���/��,/��+f�f��e�E��U"N��7��:A�����++i�Ke%H�5:j���؟��\�d�:�d]�
�y�8�J���F�@���D`U�}����F�F����X1�����d6�4FXǗ�j���6�4��ѧ���bL/��şg[!��$5r�[>�=�O)�˘q���P�:�&x�=S�@[�z����?ijS+��-���7��w���w�-�j��-�����l�U����_�nX"����IͧW�����V�������&#��Aba�i��ݼ�Ky�޿��x�C�����ۻb�[���1�7o��9�\��vr�ٝ�|�o��SH� ��Wd��~>���e�W�#C$In���R���O�wN�:;�>��0�������N�>X=}s���ㄫ���	c&���I�������^`�C��Âj%��'X+��6q�=��/���Z̆C�6Ɲ�1�ݪ4���*�bga4�)@R->	�kUp����L˹
vQf����W|~%�i��R�S�mt��l�<�������P�f�[@�j�;��-Z9�A�f�~7e*��%}8�O�T�zN%�k�u?��������ea�U._��6��_�EeH_t%�݉��%���r��&r%��G�uB��c�e��דS[�%�s�2�5���W��nϫ�
gjȂ�x��v໣�Ux�x�*.D�k�S�*���RB�]o ����w��4�/�X\ᶦ�nO��&�D۰��Ե�x����B�D3��"�N�ߌ*�)��)��D$MP��g�~�'M�dF�Z�	K���K�{�N5�49X�ϺY��d����Z��p�6w�v/2jES�258�Z�K�qQ8��h/��%-��7��f�şr�h�!��������1$�پ�1�'��
0o�}�2�QI�);��ֲflX�4��L�\��:˞��T�&0:��?�Ƿ�Y���Jۡ��^��^��X���$�����F���?X!�VU�;��զO��n;��!8Y���Y �Q(Q���"}�����y��n@5��g#��C�fA	�\.͖ۗ���g��'K����e0B͑T�@��]���r�Ǧ��:[���CA 8pG�8=�gA�m�@p�T��j�fQ�f� @u^����O�O�����A]7�c֯����n(F�}d�"ʷ���V���,Q̍\sU���u�bw��`_M�gy�,w�F᫏�SN���h7tT�t����n�4����N�9�xȏ ��J������W�n֭��bJl%�=�*�,�́8ժuEĻ�S.��@��F�8ˡ��6��Es���<�L;nk�o8`,���SM ���0ߗ�.\k�b$ʗ�Qx�Z����0uڐ�,����U�f�I�!�r)�QVl�.F��Z�*�w��^ƥt��by�s8*}L��4���l,N�+o7�����X~��Z[���뗫�Pn���MݿX�h0xq���\��Ŋ�(��m+��6 V��K¯j�Q������|hh�)�s'���^ˤTI�^����Z�D����0'��K�X��$ԧŲ`��^I�J�:���!��v�U�&����jԃ�o�u$�Y�syK��-����{
c�%P�9��r�hDP��� ��*��`v�N}���3�kEHt�T��<޼�F�W��R��k��~i���j�����`��ߎ.�$|HD���߀�ߠ���@��L֦���ӳ�=�����?S��rL5b�:^3Ծp|�al7�[/��yx� Hb_���@]	x��9�˸��fߔ�c9&�x�6���d�X�y ��?dI����]FQsu���U�;e�i��vL ��G��j|���M܂����,s�������݁����P_�|uR����ϚD�5Ϛ��<#�,َ�3?�#d�<d~��Ɔ��8�W�k��!��9���fy����Y��R2�kb�ó�Aw����b����vK
�v՜5�~Fޕ����
��b-��>�h�[�g����-�F����@�}N>�Wc�����!�IuRwP�:2�����C�S��TĚ<���΃�s��W4�t@P����c����p`�GŃ�Qo��W������C���KM�ձ��XĖ0�2�ؽ�@Xϥ$c�-ӧ���N��]bA����/{Q�̾-�k�,̌�yXg��k�Mh06n�I��x�P���_rcY����jb=������\r�iF�p�˽�~̞t%�n��>�mĒ�U�:���|&�3�h<q*�Gk�U��>OF���D��rNK�lǏ�6A�Eβ�4]�<q�͞�H�-�`�I�}ά���_�NW� "���������u�3�����Ψj�7�{{�ݪ�PS������L�ZW�(�9�Ί��gw�Cϊ!傭5�msn�>�:o��'��W>���