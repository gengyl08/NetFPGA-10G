XlxV64EB    244f     b40�3��9�� �����|�0���#�}��ɣU�1��E���תdu�L&�|׃�B�%��J�^c��b$-��3l�pێq��1ɬ���x�M��)�B�<�q���p�吾'�5!T؋�-��F"�{3�fg�@g�S���ծ ��Y�V)��d?
��PRDLX9�A���]� ȭ3>RO���U��7��Q�k?<�+�;�K����~�����:h��������	��)]�AK)hc]J�|��W��`/yj�d;y)����B_��چ�/���1�����qRu��z����2�耕�ݲmY�vQJ\���3������� �V-�^5*��ꕎ�F׀�( �"W�BWz/�ݤ`�9���E1���O�v�'������7dX�����a���		��1��k�0����lX� �˴���ց�H/ ���
�����9QO����A�����&V�+ds��>].�3���"���}�O ZTo����
;T�a�z�NF� ]h� �PmN���jR���S�@��T���w泇4�%N��r�1&n�Dv2~i�͙>�Ng�Hg�"´���ÍB��;O'�l���YY�>�V%�[�;��M)e�zE"��?FO���y�<�� dnl���� !"�cj
\����t0\2��GE�`����^��[?.=x���y��B��(�J���*�����@x�#x��N�j�)�p,4��Z���y#�{�����k���G�q�riN�17� w]��78�b��2�-�0���O�����
b��5@v~6`�t��e�
_,X&H���:�]@(�2r2&;w�QX�RcUB�!�y��#lǚ�����m |�:}����Ny���&b򥹃�`�&�^ C-�J�˘m���L�����$ٙ�ր�ЦGrYmU%��U*�v��M\��d�iW*�ym��Br���?��	
lM�H:�����-�G�('|�r,T�����(Α�h���RĦ�9�
��dKH	�u���d�,ˠy�u��7�����V�x�ap��8��'�8d�6��1:L�;�8�r��4�==X��?ݺ��֟�y5v3��ڂ��� �L�I/M�L�l>S!��M�^ڐ�>c�����F"¡v ���H��4�6��8yn�ey-�'Z�o��_=�s��4�H�c�a	x�O��[υ<�Ͷh�w
D5+ݢ�㿃 or.�3�V���Ӂ�9��f|0�w=�̇���*�S��8"*��L��T-�W��y��a��>~��ַ�V��ՑQ����d��2�}���<���C�A�Н_J8�@�4�ɭ�^�#��N�Ͷ�5�C���5�_F��r���<t�yB~�G:L��U��]J�4����)8�fJ@��ڳʱ�.�x2/J&@��e���E�d��({_I?D1*N@���~a�/n�P�y�$��dӱ�5�����+�_BC���c��1�G��+ ٿf��_^�Ud�E�0|H��SC���"Op�	�%���=�(�[��HX
��\z<1��p��ֲ�{Е#�Ҿ�)�L�n�������qiHH�R�Ӏm�ڹ}���� Dh�:�Gc�ɶ������T;��D��~���O��,r)ߜ�2�e�b�fT�������ٗm ��VC+�ꖻ��&V�,FǨ��� f���"f|-����,��B���4,������d�П�mF3�C�_�����x%�^��d�^����BE���+����~�^��b���3b�"���Б.�Y`�Ϗɪ���j�GAhf�H���F��R�rt|U��:� ǿ?�mc1������QU�V�hb�<Lw��oɫ0Y���:�0WPXf �u�o�+n��9��:���������&ʖ��z��N
2d�&GzIt�9�#�Y�&\���ø�EON@s��(����,���&��y�x:%��@�XN6�e�������1��V��?ud�S�oz�b��9rt�$$�B���'K9����Wl�?-؀pu[�"��}n����V�'�j��}�t�����,.)L�AU��m��؍�],d�\�P���WH���j+)sT�δ�+k3"�Y0���H#�8�"��7~�]1~�:��(�|REy�H
�����v쾎�6�LOh�Du:e���[��>i�w��ꅤ5�����2 ���2[���y��s]Z���})�$����S��`}?$5!���x�?���pV#���g���51�Z�l�-ܤ��D�H(_�+�1�ƨ�oH,��N�6��F�x̒��a��.&� �҃�Y��@��m�~���ˎ��W�${�O�r��Ō�7)x�4+
q�`E�N���X�4=�Lܘ	AN�=r����,�R��`��}�?��� ��a�Ϲ��+�+	��b��@��@�`a��y~���t��z�.�?��z��y��):)>P��V��Q����-�$�u{?�g�p0��s�����}uM����Q���s�"0{�V�&a�s	�`ܑ�\��w@���8��0����!d!P�e�(XE�+x�6y�Ö��{�j��5�Ό�x�Z�N{���5�UtE����V��Ŗ��ZH�P���?2�!4����O>z��ڪ�B�"���� �a��3v��v����U�\t�O��"�3���R��k
�:�[����X�����<��f���ʠ��
;����#�٣����B��j��|�m����H4�m��"�rS���>M�Z�9[yn���g�2�_�F0̀H{�$Ő�ϫǢ����L��ܑ�(����������