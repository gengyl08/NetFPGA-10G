XlxV64EB    1871     8d0����L@��k�9�3��'#Ƃ9�hμ�g�k�w�ɨB5j��!��V]����6�Y&0�܃鉮]e��7���~�K��N��jn~���탉��˘�)��$��i�%Ͳ�V��Y"��J�{�Q���Y4���0���v
�2Qp'j��]�4W�S>[̼�"s7-=�)�ƛ���ٸc�r�qE�����D�W�3�D���v{n�h>�:}�����A�_m^ � ��}w�ZI���e���tY������>�w�R�rM�_F��jE7.ň�?��ɋ�J�$8���5�D5�q��Ry���^a��^=��#X�:��J�,v���X�Bo���4��=�y���vkr���������&�PC�zx��f��\]�(
�Ȕ��1s�ɢ�[��W�$ΠFG1"�)ʃ�U�[�s�pD�%2����
#��8c��ݨl���{J��Aܔ���.��-��	���(o>��?b���-�ښ��/6z�<V���ꨵ�z��Z��h�:/
���K����@)hK���(�-7w6�V���s���f��d��S�:�+.��1��Z|�f�"'�OzۡD�up+V@4F��n��̏�:�H�HI�H����|�]>����P��GR���0�/�G�x�W_�B\�H���Fy4���i��*� ���ܑۨ�^M�!J���B�Qfi���'�9�u`�͌�:�B�ͽ�i�a�f��14s��Y�YЭz p�u��k~�@��7��Ky�9���C��^�Ҹ���n��H66Q����s�6YE�$�#b�r��;d�|�q���On��&F��L:����<ٛT���/Z�ؼ��u�M��w$�������M�ɰS�DނW���o�mu7��Uپ��I\�Z9���Jg�@��0p;�MW�#�I�kye4ذ�$�=%5_�_ѳ%�h�gÃ7��oM*�'��%�L�m��o�<�7���:�́鯿&!yc(��k��r��8�� 2���_�%����ޛ���E���jT�B�`���0h�^�0/�6��bդ�)�F]~tƾ�m+��W�o���P�Y�+^���G�t�Ӎ�d��Oa}����C��ݚD�1l�l�j���q�,�TX�ة����}|8qxjc�' �$�`��!����I_&4��k��~���g��{Q$�Wm"f�z	��JHh�H��~f'��qmaV�������'"�è�"�B2a�������a�)��e��/�����@<Q=YB�����=E���J�]�ݍ���� E��$����Z1�/j�!)x����s�9�Ww�CPYu���#nu�J��=d���۶��lkzm��M�0{��VӻeZ0�Y��c�<|�ς��d�
)b�M��,&���n�.y�}|9��:���ڬ��.�^&*'�oL�}L�eY�s.�$X�<�aT���o�)>BL36�v�B}z�]$�|�n�*4V��4rW �_Y����k����`J�;)�Trp�;7�H���j�z�KO�N5�L�j�b�5U	��<1̌�����1�|P�k��}�\NH3��-=�?}�d<���0V��b�%���Hqz�t[ÿ��tU�У����eܱ����{�W��JG4�M����1"]qֳ4D� ��>ò,9����f~�6u(�׻џO��-���L�fѡ�b��:���Ur�����rtx�*f�k�����!�®ﱀ>��[}��Jk�(�Mt}�m�UK��,V��M7�1n�*jU�� �װ ���S�P���ג%���ª�lL�'�����Z�1�H+�хgǔs���E�~�s|Z�@�|A�j.��)���K����k��B�MsU��$��׍��WD��@�Sk���~UX(��!�`�Q��!@!���"i��jzP�H� aз�������	����aյȨ�3_�b
���E�1�ĚQ��_C���"	)�]��q���t5.�js��-h��:��?���G!�?�IjI���3���=� b�,D?^��(XX�@��� HD[1����/��yL}�������]�' 	������ [ۆ���C9�Q�E2/e���u	*,���ٯ�2~c�0no�߶й��#j�u&:V$&��9�7�_VŃc�Y-c�r�3-O �<A`�k���)%��C���ӻp�T�Ǎ�)p5����'�ǤR5 ^�c���Jt-Mm8O�	