XlxV64EB    182e     880ft�I1��|��c�����no	PA,��@������ �A�f�m�E������2�K��{g���Wn���e8��Gڭ�	���L��/���'Y�l\R����>��8�J�᣽�Ԉ�����-f!���=���m����
u{#��dB����� $e)��p�R�Z͐Ґr�W݃]@�I�0�K���]X��F:���(�;sF5	h#~#W�uӅ�Ǣ&�Á�<%$�N{��&�P�#���&�I��|%E�TW�$�
���HE���ں7=�D�ӕs�7�?� �l����f̷�xAR���Z.�^�D����a:�Y��/�n�8�Ӫ+��2یo����.濃�G*^��DXP���N�P�� �-^W7⿮'1)���-�����]��A�UҾ�!�r.����h��R�>i��sݴŐ�x��x��|����A��lLbR���',3{e� I�w�g��
D+�~���������_��9��24=Ĕ��U���]�c�4��R�DӬ��|;=a'�2L�e�;�}����c	y�������=uJ���F���*��3y� i���(��H��D�r�!9��& &L����a/L�u�޳Y-��_�|s�
�6
�4(j)�J��.s������,��aֿ}@��4�~�	�� 1�&JB���?C>"���Q��J����O�A�%��8����FL��+��L����؊�d��7Ё
��2�l%8���$�*�
%
���p���jN� ��e�P�	��R!!�~�C�a=u��i=Z��EJ,?��ʧ��_'`��;�����@]�֒zC,=��zݥ�TUpk��Ya�;��o碹%�c�.~��d��SUA
.�c�Gf��Pf��::?�o9�YD��:A���Mi��p�� �-�����<ө��td�/�S�CM���N����[��4x�`�,]�v@�h$�Gu�"�	�g�B���b����h�U0��	Y<�����!8l��ej����@.5�ai4��M���6�h�b��22�&�]��z}�1�_�E�d_�V-Ϙ����������h��r���>U`�y������M,�/���r��xo��g��f�{W�뮯��*K*�}�y�J���5�/59�����u
��S/���VpU�@IU��`V)�Uڬ���mS�=hyt<�9:%��.�{�jt��H�� �h	��f[&���7da<��b�A�	5A�8���ـH�ڞv	��!G];�rN��c�ilN ��� Zm�� �3v��D�u�,i|�0Kc��
�IÑA�6EJ��Ӌ���Mu"93���{0x'�$���c��/jRO
�'G�R��7L�y�x�U(�.x��CS ��Nhv�����L)�� ��H٤�7�7�@WZF���6�I����Њ�	�7�swBRB�`=N���j썅B��*��\����Vp����X�"��1�}�X����l�N�(�rnP�!�3�.P�S����>L��x����}�CQ%���f �XоV�w���,�+��X��Dm�N�ű�m�y�V�~E��hUz���������Ԏw���g=|$n	\?�⸈>�2�q񔈗�5i^��)D�|��3)���d'eg0���,�v@v�� �����m��	�x���A#- [N��Hf9.��T�{�:T������v0�c���[UZ������[Q�
�!��4n|��V�݂	_"^O��*���R�ek�%�v��1.�q�=�-�`�j%t�[���c#ץ�=�I��������\�����Ț���_���FU=�x�ߏ�7�obe��sv�FsAiyt)}��C�`�j�c�]|H��Z���?4)(
#Q#����\հe�ޓ���֋�s�P�m}�~���1h�od�afu'ג�=�2�r� �:Q̌��J�B�d�LN�u���uP��?sw�Fym��w�u�����*M���M�'��"3�O��цf�g�Bjn	ú�P1H�p2OM#3u$�b�d\U56�DIDx?��,�"`��!����C:��m��?X\�'D��%LD�(ӻ���-�<&�`�À
' ��*6�۲�@�����T	�2/$��OZ�vX�r�Z.�H�y>ԩ�{�è2���<?���