XlxV64EB    1e37     a80��a'�"_�j	�m��,����`]���QQ���U�%�2v�]HƇ��;���YX���l�v|gt�OF,�`��T!����r'upV
�䒰GeN�b����iM���OHm{�=:�y2�kg���o���{+��0t�ݭ@��[���p��c���>��]�3����M��OZJ�h����A��������prq��y/M���Si^H�8�e����]m���2�q���{�sʐg��띁�̘f7�a7�����x�g7QfmlE��H�����Wjl�Щ�m�=Gc��Ι�@*��<jDi{�5^��fM9bV���Z�~h��h�\y��N��e�cG��}H#�sx�8�:& t5�"s'�l����;�����<"d� ё&��O�B�ގ~\?���P_�$|S�� M)����X��!"oӸ5_�6��U"/��_��l��j��<ׁ�8�9cҡR�,��V��h�EK�fD�FnI�fOb4���I4M��,t��Y@���J�FY��@��5�'���=�E1�Av6O�O�]�z<��B�������li^}��KY'bP�q�^^��?��?�䀀@��ܯ[;WG@��xp:]W��&&o�Sn|"���&x$F7c֓xN@p��!�\x$����V����ԣvR��PSjE���Ε�}�.6 �,�5,I� >L�����U�ޡ|$�PDf�&/&.�����5٨~�)�C���\���>�b^�������=˃�ù4=b�B�e#3���v֢%V��/�떩S�����Y��YTD5|��t���E���B�-�ǹ@�e��CJ򍔀@"�8��g��hi����1? �UqP�k�u�z ��x�0�����ڷe��1�F�s}�X��X5c�.?(b����]s�:A!��]gm*�:'�ъ@��hL� mF�i^�I��컡@��`�/�ӧNA=����K����V���V���]���g��^X[f�D�A�7��X#�}�p�om����&Nh&5�,����˓�{�*X��� Ke��3/Z�z�(�u+_��8�өpi\�n��
�WTYe����OG$<�/{x>_B��窷��x�����~
:�j(��@�T���,(�P�T����7N;~f�zRPÛ
���T��	~���G�T�dG���� �����$D~M�!O@"W�~�*.�zhW0�fb������N�e,1��Kk��q����Ђ�)E�י�sN9b�a���E�JL�?5|�F���3y�qϺI/�w���>�'���V���m�b։Ǽ"^�M�-�Ϋ��O�O�"X$��|9�4L8p����J�ni��n<���E�?�Y��DU��$Jօ����LW�d�࿼��Bx�aK煎�^vlj"��Y�#~�G��%6D�a�g\sa��(�他b�6�%;�ȃ���J��?��3l81L�� WΪQ��{���D����0Ԡ-̡F�ѓ�Yt�!O9�g�Fk�H瞶g&��Y��\\�By�� Cm'��@�o�4?�yH<��JY(ϓ*)� t�2f���%��� _"�|�o��B�y:���B���z�O-��Z�0���F؄�:i �ڭ���8�?z�}����)���}i<�IҜV�r��֓T7������l�ި(e�Ҟ�󖦋*__���َ�+������I����f��	G�)@�����*��XeFT��Hu�E�#B�|���Fk>`� Et��}l�-Gb;��y0�C����_~��VY�q/n# ,!Y��ČT�5~����"��Og���B����ky�f���ޭ��������3���j�p�v��tmv�s,M���)RH�;s����(Q�����ڠ�M5�ڤ4�w��?�ذ�;�k>�UD�7���3������/�̊ǦZ�B@��<�Tø햌��'C�+|]�p f0�iv/�ka�@�Ri+�G�����K��Cc�B���'3�|���OP� �8b��m8>�G�9��Pj����0/�=��X_5�3��}8�g�0D��U������k��@넚	��]�-Îe;��\���P�$�{���(�����L�.)��k�8��ݨ�A�W���:� J�H�����-%ď��F6lVLћ�^���y��ɸ�\4�W�,x�a�Z�)��rkx�"�i�rJȤ�P���g��᱄%j

�	r�`�*��+��	5��Fw��Y�a�a������g�i(����a�p�RV�w�,Ś3�A�x�f�v'-���?i$�Μ0�G�b8⡄����+�w;HSR����o��G\k�C����
�V8yvj��f6�@���Z��� �,��Z�Rddێ��=�	P�4�4J����O#8��!0T��b��z�ÿ���G�B�C�k���� ��@�����+�[1с"4�I���\�PfG/�%������\����U��Ӳ�_�ji>o��IY���m��!�.5�a�����@3� ���90�k�$K�qZ�!@NC��V�Z5� ��%�yñ��D�J3T�%+W��``p[���'J�5��y(l�{hq�~�����{*k�ၓ~@�pa�g�#���_�č�B�gz�ޏ<�id���6����Y��%c z