XlxV64EB    fa00    2fe0] ęB��&\d�O��g�Uip\�r��^��j�*�䀸#�2�y~�6ҥN����g ^�l7G�n���������ڠ�u�x�����w47!U�0bU��'Zx笲�\�.w�8�D��'�������<}Yy�N��ㆥ�����]�jm�����B��'z�Y��ppM(ol�C'��(�zD�q�
�߻	"T{�ܻ�?�ݗ#��4�^Ucmt^F��.��$�������I%�<?Sq����O_q8p��y�'f̮���-��ִ͊O����h�~h����������W9���HVT�퐖c�?�_H3&tOqSd-�{�Po�"���5|1(�����9��D�=�{��~$Zt.^Sp$���l��[5�p&��Dd2�i�qE��hT���{u&���T�b?]d�cx��
��=���z�Kd^�_N�{X�)�8g�P�V��g��b�ä�R����f��52���~����XdGַ��cS�����N��n�_Y��gz������n��:�0Y�N#�2#)�I5���z�?�nu��������r�ZD��9\��=xX-ik��а6���l��=��	��Ϻ�Y�Yұ�I�A=�SZ���vsMK4ae���@�B0W�,�	��Z�i�Tn	�@:�h�C\�}����Q��~���	�T/W�&#8�kM�S��������؞Ι��
Ƌ��@�!���..��W8��(���}Lg�SLoo�1����n{N�Ax�a����Σ<�ʇv����[�+��B�(�~o��+ܻ*��?�}4HͼA�q)(C%�������gͺ7V��j���qk7M���z	^��_��o����ܮT�`��s�k-�I��$g<̃5k����`�hA��}�'�3F��`�G��տ.Et�e�g1N�"W��5e�=ݏ�'@�j�CT x|g��3�:(����iU�Ř�\�}9�G�>rr��������μ��k��.>9��Ɲ����V���J�`��c�炚n���L%&�H~K'j?��pM���^AK�/���p3�>OTd���s���~�4�BA�*�ILR�����0A5}��m��ζ��5@�r�a�8*I��o����mkY�?]f.��hqw;"��o�h���~2��JaYFğ̽�~��}=�=��]��M�5���'�rhߨ���2�$��h_�q�tM����J2�Hh��ع~$-��@�T�����N���ˬ���Z���
��>�*�mĝq������~��1�^�b���eπ힂!�4�qp�4M������DrB��<?��_�]Ɔ��T��|p۽1n��}�%��M��%����rڤ�9aLi�C�v�0���T�"�٧d����騡[��J�\��x�҃�*2�n#��� e�6V(F�Do��M�+��7�U�j�z�#V��EU�%<��Ǽf1�_Z�Y�.2�|�Z�W~����,���M�9��ą�ў��k���.���xH+��4 �K
M�E�}z��fI�x�}�6q*e���P�\{��[&epεqI/� ��'S��&0%C���O�b��GZ2��|�}|v�Ɓ�Dt�~l����\rmx�;�R?�辣�`�|��+ݾX|�)L��3Q�ܤ7<5�;�0�l�:�G~5ؙca�l:`R{\��k��m�0�)CQ?_�?�PGIN���0
j"�Gc��.�����l�b�既/i�`��~=f6������X'�i�;���-Fa�{��ю��\<,�7|�	l�{/�۵��1���Uτ��J[p= �u��T�����;IrFDt ���[6�՝��;(��qY�x�RԢ�	'�!�ddb����\"\�(�N�\��^	m�=�؂�>�?�r� �@�:��A�#���c��o��pN*؋�*�L�75��?�~���Sh�k�:hd�k��e@�y�փ?�ix������ʟ��ʴ�p<RQА)#&D]���ϡ�6F/��t�B(����iG ��g���T��k쾐����=Ġ-� ��[C�Hy�8/�_���&ٮ;��&=��f�Ʉmx��6�?�X]Z�V YT{�pK��*>���AGa$@D���2��so��J�`�n��Xݰ�����p|��'�d����Au�V�{�mu6@����\�H)�tʖ�=�7��@�����)$�Q�Yٶ�)��/ǻ�V~^��#F;7$XYp��"�����B�a�?�P;�:=D�)�r���eÅ8�"�(�m��Y����X��OP-KZh3;
�X��/�!v�OD���K�&V���RUFFAs�F^��m* I9/BY���ч~3�WN�;t��b��)K�^������좋
?�;���WY7� qR��V�`�{��-c����[�ĵB{<�	�:t��1��'V��:��+�	HՏ=*��1��H���.c���%#� m�E�d*��L��,�&�����J�Sm�0;�fX������ P0�&M�ww`'�m�4�P����F}!�Mm�S�t��e��,��R�$s�oS�
�*��-�?��6njH�N�T$%���Os_�������BD�V�I�>��<�}�9y]�&F@�iCC�N~j������wM�R.��]���13HgG��%�FA�G�'Jw3b�%��4��"�t�����I	�M��9[&9�.`�/��,���-��'�,:�WiI�I�f����i��;9gf�V�h�3zo ������w����=�"�ڑ�_�*��:��oA����I���:l��ߗ�5=�C��v�4�GP��6S�*�:���"1ɗ�C�pe�%CE����,cEox���g�|�US7����E7�0Q'�/*Q�BZ�g ������ʷ��]����E��>��D��g/oc�W�܁��ӿ��R6ݿ�AX�-�t�2�B`ʃd���6�Wg�P@bԎҊaU���ƅO�<WlT�fэ����8�h���^�v1oL��������9 �@H��'���SėX>/��F����"62�]�!1��P���p4�je���gP��Y}A쫷�zonM��0�y���������˶��Q��«=��ֵ�S��Yc5>m�_9�[P~oo���b���e�#�2�����t?�$�0�M�K�
'�ƃ�7�,9 Q�#h!i�ߦ��5,�)B���K�b�$�8:��'����W��SF�FT@J�?Oo�ӹY��D�F���܇ې�����Km+��ީ^���lw�9=�O��O;^�m}���C�v* ���\�t�++&���(��M������3L/$���=���-Z�Ž� ��(��l��(��Ķ��[��J:_s�}]�������P��ov?9�|�up,�[xj0P~m��L�^`�.+�Gh�����	�S���E�r��z��v�)`$y=&acԌc`�hQP�j�/`�QY��w��]�Dvh��y���[��s�Qp�b��mg&9��V�B{�W�~��%+� ��"����Vm��0�	���&��H��J\���������t�0�Žo�� A���9�X?R���Kݤxa�Z'�q��bN�� (�M�'�߹,Dp� ���
!���a
=�1��,{�hod�甀�Ux�z���cP���*9�z#�9�~ !������;J}n�/������������9����yݳ	-������f��p4����maۏ��?�aKT��5YDQl,ۨƼ�)ӪQ���i���R���ߏꒉ�~�#N�[A&�_*�*��lv#�*�ὶ$�eI����a�tizI��U���~vȖ������u�Tl]:[�w���1��IMh=X5!�_р��>��ƽ���a��0���tclE����F��Of�j|��#@4_�������ڇd1�خsf�i�����?�6?_!�c�׽�b�3��3?ċ�m����T�����)��������DV���J=1����tN)(���������%��+Z�ڃ!�7��;��O�+2
r�afG����Z�����1�v]%�?3S	3"ji���L�O����2B��8�A�e'"���8��n����$^��9v'He��3��Pn͕Πr^[��(O�s}���
���l^"�����]T�x}�0bf�I�.#���8�pb�Nd�J9�(�2Ǎ��AE�B�㑙c�lE��K4�.Mq)�����ѾI,�"�8E���tL��A�����<��P�S�_�l���y�Ȅ��33J�~�񗚫�ط]��!��i��]%^�z��V+�A��%����w(�jdD�A
��eF���N�y��j8o�E��!Y^��R�d��1�J�=\�bw_�.��%�9��,¨��a�Xx|��a蘧�Yl	3���A'
o{9�����RR1�Ъ��2�(���[fa�㔑�	$E��,�/p�Ѵzy�|�����`���(�c'�銧�R��:����F<)
1W:s��=�`��7��"'g
�L�(��BN]���1�6#�B���E��������NrF
����N�)۠��Wd[�+5�?�O�k3@O��� nK~�z��]5a�ėS�s�FR�`.V__X�8S:���
��Z�0�6[�ޚ����!��>�y,~�ukQ�O�x0����uGB��n�T���}�������x2�A��2�$j�WL��W.l(�t�#��-9S�*K�kD/0���Ώ0M�ɽ� ס�TҮ�^8��_)o�5��Zvl�x�Yu`Q�~�9��˒?+g���F$�јm��(�"u$o%'^h���gQN�E�Ԇ�@G��?)��)�iW��w�t�Y*.OJ��D�L�p�պ�:��K����m���օq#6A����ꩣ�580�������O�%H5q�\bHl�X��Q�K!ݠ~�lȑ�*!Ű	�%p�]u���*�"��3l�]��~w���$c���4��B�gg�AF���o��&��'F��p�Օa Pv}�k;]l��!(
�i�}m��앶�)u�E&ʉc˄ y���1�(���Zݓn¦[d���tͪ�)���(f��ژ�|0I�[�a�G��{f!k����O B�S*����rV�qȻ��]ͤ�Q逞���&��r��W�3e%�)����j�K[�>N6����̓�֠��K�ҳ�=����.Y9�����r_�SX9�~_�GL��^p�ymV�T�仗"�[R��O�xCw�����Ǭ;�de��`�<pn����8�]�j�,�/�x�w��;�FG�PX�ʤ�u�y�F�~���C��l�b���|\�8��� ���C�#�1���,��f����*�D� 5�0U]}A�$�*ė�|�$rΙCtG�54�al,?L���u��p��)qsCsO�gD�ֹ��&���_B�VEH~��)���<Yǩs����7�wN7ğ�x���<��z�d�w+4X=�C���͆	��#�ϝ�հ�S'Dذ+�N�L���6�TvU��Nh�(]�1�
�TPj����/.��V����{
/���6�j�SZЀ��T޵�wRIz�R�>�k]-z��|w��X�+J?n?=��I��D�a�Vt��@�����y��^�&;�Jܚ1���B�˗�Y�� ��=���k�|K���n
�\�>ܟd�[	*i�Ҵ����{�I�P�4���1Țgf�I�_dW���;$e���9�
,��*���91>�b�W�V��Q���0�٥71Q������jd��ŧ�q�N ���e������|��!��Gt'O�Rh�?y'\�Ï��cQ��w��=��̰�����e[�S���[��[Q1�p\���)p�����A]|[�@a�ۊF�����)�B~�����M�&��Up��B���ф �I5��
�<�G0�b��0鏂��@��7���X�y�p��{f�Q�	6s�j��Xǣ��<^=\�����<�!�nqx����1�F9㫍�D�����"��2�6���4Ҍ�c�(-�6&Ċ�_'�j���5��؃�C�y,�������orE,��t�ȹ��.����|�-�*Ӟ�*^9��q�b��Z����W��01(F��N!�f�y�PM����n<MtQ::P�3
W0�*��#�{Y�����B�k����Q����!{F�F�h�i���G�j�ច'T�  ,��xtjЄ��!�L�����;X/F�E�P������Wd^�f3�I1�|Dw&�0`��xh�[tN=ai֫������k�1��������U�ֿl�,���ŗ�[�&�m�4��g?ڤ������@�7��#�d��̒�Ť��T$K�~�u�Y�������ۄ�.�~I�)��G��pã�t�7̈�X�'A�-z ��a�Lva#�qp����]�X������\�X%��Lx:s��W�;��vMZ�5����U7;�d����F&�*Z@,�oD��S{!��_'"5������`��,���7|��D8'����J4_~�O��\���k�&���.R�� �\�ɉ�i�L[���'7�~O�\�s� š-u0��ܡ���˿��+"
w��9kT�ӄ$$D��CMR�{+
�G��<}�TBr
l�E8�Q�D���0���a��>4��Ւŷ�a��ݼeP�K�W3XM��#����r!���d�,��k�=b$ו#��rwUA�[�`֖"ٓac36������^#�&��6�'�6�^�! (=�E�8A�וֹ�oQ�Dˇ3ِ�}Y�������<rܣ�)��ԫ���VQ������<@n���sZ��Mvm������nXl�p��1��F �f��K�c"f�f~�&~�*�I���gO�U�	��[~=g�Z|Cu�b�x�e��B~�1�uQ^[�cv*���?��{^E�S��)����#=�7W���m�k5�����gs���8�S��jX��e���e�o-��cc�l
_�ɀ�	�$��vH���ȧ� 	y�,�ᪧ̔ˌ:FbE�!�􃭏���)U@��-���ә_c���Jk�g��In���s�P����;��G/�;�i"��ŝ�/�|��2��;W�~Oy̮ї�X�+��z���#��PF���.!Z�¤�P���E2����чz���0�]���T8m�����a�wJ__
<2�7�|�B�)i��ɵz��&z�̓J���CL���}a� �Yz^g�ۀ����>�m��u9�Wi)6��˂~��W5��C�76�F���B��(��'*qg��y��~]��aV�3�[��Un~�3���Z���;&��������<e�����p٭1L�t��6�Pn���K�H4����<�V�U���`f��Ԁ����!�R�¢ �פR=F�r�2K����8�F/\�j�Hl��I���~e���+u� ����Ԡx�~[�s� �δ0�с���R�>lw*y��U�yӭ?�y�]8��Dt�sw�a�HI��	�lct?&�Pe�>jn~����� ��^���CV�"�
����#�ƈCm��X6�{�W� ,W�*.+c�����)��5�+d��
�&�{����0�.��/gѪ{Hά��U�ڏ���OH�����Q�DP/Mm�µ��+�����n��v��-5B�^x+TG��5�5� �|sq�.[I	���K�UB��ٸM`^EX�(��#C����]pi�Fҹ���y��K͜R��I�~y���\���`�W*?���+f�9NIK�P3�R�-Н��Gҡ�/f�ե��D�+(n����ˣD��Vgi��U&Gd2��=���P#I�6�z\��?�h�C��!�Gĵг:�м�q
���B'e�-��Z�L���F�+z���E��$��l+6�e�)����۪��8[�(4$�݇��
�Q�y�����j�N����):U�o�EZ��}o�f_acTq�1���Bn3�GΦ�%�k��!�c�{�.�����67��̲��X����(;[�yxA[��J��Uex<��-�C9�@SD����7l���.��Zڎݞ��Q�"/�CW�#��g}��"����r�����(Ea'�@:p�!�V�*�P�7�����d�m��t���{�bT6עk9�9vrAg�!����٘:��.��z#����%{��y�8eΧ��6e���7~��F��Q��;zjCj��XXt�ߥ�|'�aV���`S��P��X'4����2> t��
��vK�;ޛdLB��s�I�tt��~I�����\s�f�����wX)���2���^m(��>��0oSP��3������qKE\��S��1p�DKKb:^S'wy�̕g���T�y���׭�8Eй0��qtuB&`e���1���f6�~�{z��+�m����{�P� ˆ!|f�W?��g�����g7">�fkYE��8��u���إs)j�'�i�I:���9�Q�sر2����7�ʄl����tT�|Ly^�5��薨���j�ucC[頵�;���ͺ
r%�mCMIv<RUs���?0�Z�S����N�����+�ȷ\J�Oey��=��A�9�!(g����t�5~ǝb�g��x��ĵ�V�}F\}c/H�Yl�9s��C @9³�V����%U�X�U"Ø��͵�N�8��E�-F4cD�!�{b�G��×�����Rg��Q�bET�JT:��n�PK!���M��B���"��M�4�w��)xڻPÙ��9���:�l[�Buk�Kb����	^#>�M���M�ó�p�}Z'ڞJ�v�O���Z �XDN��b+7�ፁHI2z��ɗ@)*����q�i�C��-�^[6BqG�}������R�L2�܁��U�N���T���kO��*����l|F����D��I���Hs�_v4ɐ(s�9i�3_=�U�<h����-4�c��d�L��ט���$��F�I@��b?bv`�Y5���{�������)����4�K����ۻ�6k�'�A���M��5���RJ�w�B9b���L��[�h��[M	D�V��(���ɯ�ď��;��:$����� 4TO\Rf����y��,�Pkܝ�h��҃�2Ei
�I)�hL��ߒP�hp6;G[��U��\D��Ml�����(�>�����f[D�4ƞ]���)��\�F��(��y�G�!/7�%�WUcpk̄�k`�j��1��LA�=+�W��%����֏���\[o(�D����~��+'R7�Sq�R�6]D�L�m�ԫ�s�e%�b��}]�t��"C����,�����tܗ�6����b����^vZ�îI����0��JU��rl�U5�����A��8Mzl��Sj�������e�����!@I�"����J3�R\�eX���1�­f1ÝZ��qʟ��ҹ@g�9ķ+W����("�!W�B��w`9|x�
�|{;R��`��N<g�~��S�{�Rw��vN���1#N�8jڲ��b�� ����M�#1��
�_ڝ#î@v�:��3���&�'Lb�E?)1�}��-o�l��SnEs1s�}�&
��Q��n�����3H�2���l��a�^�~(_��3��K��w��;�������+ϵұ��OY��2A�����)7E�Z>Ԫ�T��יo1��W�w����QpQkh�Z����P��Қ�	��	�ٱ�g�ڂ�L� ��@���m��,*LFr���%����Ѽ�
xy��zZ{��zgt��Ëp��U]���y�c�����h���kr��w�z�Y�����	Ѹ���;(Z�� �o�>�I����V���ހ2Ӽ-�J�`��%8���"y��ղM��#a�Z�8ώW�}����p�Y쬡�>C/A}����)�	&�z	 �ё8�>FM�]VB%�7�dp�b�]O���H�X/#[�?�_D/C�FF���`č��"�_o�ا�c��[�<��($��5�ǰʄ#`̍��n��q;`%�W�HԂ��7��?h��{��OvP������J�*[f�5|�$<T��}E�6��l�#a�.�86Y<Zd�ఋ*���fe0G�i����b�d��7$�F�׳�3�˥N0A�-��w��H��(��::i�s�	�O�R�
�@F���+CV�p�ǿ���98R����87��w��Cۋ�N/�� ��D�(s����7����+��d�Dy�S���wR&�?�bw�F'��9tT�(Q���a7Z
�R!���6N R궁b���R
?o����l�El>P�7Y�i:HX	G�h�9�T3;�v��=m�66E��T�VbdC.���ŋ�4pΣ5�!;�_+T�O�3�]e��i���X�r�o-�G��[4��(}��?�	  �C�|�1� s�R��v��J�P*�b�(\"��)��<1؟�E�k++_�
.>���Ӽyz���������������[^V���+��t�6�6o�9�6���ٻ� �<n�x�f�#�Ƙ�<�&>�2e���?�"�ՙ�V`L���_� ��Q������*�嚨�`�ɐ䁥�k���'���U�\������{]H����s
�9�e;�?HUr�k���U�����UV8���V�����xf�o�@�7��~�R��i�]�|2K�!�B}�KMZ�>6�� � �nm��_�#4���{�Mq��F�ǩ�_�HW��I�qL�U��=��-$���{�R_M%�#8/o�D�i�9�R���9�
��j�5�gs�(��n��C�"���rϬ+��5�J������Dx�\�=�oc�u�s�o/k�F��!ʩh'�~�/@����� �d^��P�/�S��e�
��=�����q��mN\�"�� ��&ГBq��zT��&2/���h8�\W�����t��+s�%&q�\��Ư�E����|��V����H�߹�(�O��<��E_���шhȵ��6�~=O~"f����/�eZ�.Gy�ZzqC��sMo�&I$�o����Q:��?J��NM�J�
�j��$���h6�0�6��퐱�==L�p3���[U����'eܘB�u�i�=� ��x���zh��.檝��
JL�͔��E���8'��ޡ���H�k$�y;:���g���t�fg��_�K/�~R����ȀH���G���q<�� �:�#�b�䰅t����q��]�K4O�V!�Ϧ�.��8:�p�I[���
p��rQ�ϻ����W��!�_'6c�\��]��MYMy�����	�}��23��=0������c�/anT�����1G�2qs+�^���+���!і�]�=��~�@�V|KԽio���kp.��)��3u�
��2�G����JLWGJ����B�/�6�i;Ճj8���j>a
 y���Z�XI�X���vzQ�ЈkE
��'e��C�N�a��\kG�� �YI@�/S0�ee�K �z'l��W境"����>�L��b�;�h9ٶ���Z_�ĭ��:���y_Hx"��׹6ن�7'N�U��k�����8> �ʩ���+��q�Cဇ�_-'��V������@i��r��q�Ύ�S0&�ύ*�I�Ҿӿ.��Qd�_h	�&���[�(���ifA1�p���!A/]���(�:j׭���:�>b�?+��e��\"���P���7ۺ{�� �)}꧅itYW�T�i/^��/̫
�L��w�&ql���X�Sz���2;�Jv0GEw��08�8,�j�1Հ�kh2�*��kڃ�0�/����S��@�1M��Z����+�e�i��6��_EhM��"2q�3/%u�qn0d�f�<�����sU�>L(.�|uj�(ǭS���0�s��0��-P_)��a�v^&�����F(�Mt�#"��Jx�0C�	%�p�s�����n;�����ɸ���T��\R0|MQ��e@�Q��q  ���	֘tw�K��i���t՗�m�]�����]%�6��B���Xd	x��g�h�*O�N	����_�HE�u��t��*/�T�Z}�� ��D'�_g�a�����-�
XlxV64EB    5f71    1450��4#��-�a	�u�{��?l�vG��G�����(����K����PᇸFƉ=�@��Γ�QY��z��Ch&8Q��,�Ph�+A��K_:���<#V�v�{�? �{
�[1�q�N��ۥ�y�!���@\�=��hS�	�ʗ��������� �~�	�)#�s�}�/x��D����􃢦�Q�t?+����ɑ+B X�I���{�U�c���C�Vڊ��<��z����vlɈ�+����e^j�7��k���	�/R�p��_�;AC�:������ӺJ����5ruX�����+�R������1��6�)t�\[��?v���l�����T�:��M{A+'�@��x7�7J��E��x����r�a>cK�;V<�?�`.���"-��Ӣ��i�j�xѯb�@����'�V�����ٲ��*ȥ�i����?q��k������FZ
��ڍ�<kF�W�@ RkT1!g�O��1}��F+���N�Z�B
�Ϣ2�9l����^%L+;bB
D��`Tjf*���7�r�l���Ӎv�{(��m5�����O ������kz��(��t�`�(ز�93����T�a�����Q�2۲�+�[��N��H.@/��1Us���� -M���fgE�u�Q�%b�-Y7��?�A�ݟ�D�w�|I�|C� �z��H@�2�X4�b�3��ب�X�r\���p��4�,��*����/<�T�-׃��	Q3��>�p5�#3��E*cfxPӘ���0i������;T����g��C�@���n��x����㠕��aL�0Q&XܑT�3}ⱻ0�JH�^���͎e���C�G24�}�إ���Li��C󝤢Q����&��nv��C2��ȠU0����&���n����eTƚ���_my����ip���=&�2�k�+�T�R%�11�9ޠQj�9�y��њ�'���Lu�,: ko*�~�a暧�طӻ鑬W�/4����vzk+�:z����nQ"$U}&������9Ӭ�7����χ�����}{@���H�m�cH�eے�3��&�(��e+Fw#J����U0�0�)E��o�e��v�-�t��'�dJ	7Ֆ�Qh�8�u���#2�$�Ł؃́Kj΂�R���=�"2�-9<��Ga������ޞ%e�����Hd9	FU���UA�s�%)�:?n��+�N��M�28s�*��<��zQ�E�[���ȩ�T3O������A�l�X&ޞ��%���4��R�=Ҍ�����T�ָ�&]Tc��j%��� lIIZ9$��Ԗ�Z��@8+G!�u�n�r-)�>^�M�wL��`#*��סt�c�CC�a�:7�{��]C����r�v"�]�p8L��ݕ��v�<���ub��;��Ǐҹ����HѦ;�_��%�@|��o��8*����Q:Z�*kGƠ��1)�����ứՑs?����r�$��'�ޖ�s|���yؕy��ƞ�~�X�V�+B�.��;i�I��=�pj�<����N��x�U�d������i�Z0َ)�<$V�x��4p�"�"E9ʐ!�)�3�ÿ�A]��4n�t���9���Q�G���v��T_���`�2��p�G�-��#>�ʸ����^��ɍ㋬
�&EOd�Uљ�x.s���t��Xn�����j��F�hg"�&���}W�2Flpٱ��Q����aݞ
��\檺���N��UoY>E�x^O(:�֙����E@�\�9,�a&�(O��Y��a� �"��]Ѱ)���ZP��ܿ�l�K� <Ddj�n6ua]5N���n��Z�9 (i�z樕:�Ғ��w�a�fB���T$g�i�Y<x� ��g�?C���n�{_���,��+~���.���}��]'��)��SLNi�g�Oo��MH��7����@��+����鶓��d��e�A�����v�^j�̎��h�����>V�Q��0��S����R��w�&F@ֈ@�V�e�����U]4�Yr����_�,0��'�d����+A�\���Q^����o��Y�aV���{Mܥ]��3h���"�&������A�1�Ϫ�� �����z��1�I6;�u�@ީC@�-�]�� .ڽ��!��:�O*"L�Wf��hϫ7�&����u���CD�J6��H��4s��E�l�����	����>ꄈ��;�A���}y�4�(��:
��a�x�v�
�>�g�Vm���D��u�P��:�|�%z����n:�9$j�i��z�,��j�����O�)Ռ��zn�[ʶ
+��4�����9��j����4X���t�v���j�tF6�N�������i��0ܔvv�@轟��$~a��rɇ�����x��Y1���ЙQ�P�0�Q�ߘ��$��NR�O���A$OҮfu�"��7���<W7�d��:�x�$`�*|ኋ�W!�#y��5q8Y��0G���k��w�Rξ:����U��d	b���hY]��3V����j��N�<�D���
�l�ss�%�ԴK���5�Z^�$;r)h3׍1�lU���ʙw����������n*ՁQ(��?PKDV�w��^j���
�f1�O>���`�$ǔ<��%�a�}[X�ڨTSIζ��=�b�Ag���8$�+��K�n-��ٍw��f�v�? pU~���-j� /"A�1jj�G�u���P!��vڸ�T/�4n@`?R�R�@R�c^D��(�w*
�{�K�a�i���3կ�@{���-�tF0�2^s׍����8�6$��u��#Z�ag��94	x5��;`D�zy0�D���2�ܛz.wx��o�H�+�;Ծ*B�E&��ݡA��0��w���T|M��b�Ln!Z͈�
^�L��4�pPAK�e�� C�QFs��
k�K��q��d�_rt���mvO#��"�d���]K����)U�m��{�ƴ�]��^۠}b�)��#������[ۺﻮ�L k}��ѳ|��������鸼v0�ZlUK���{ذ�&�!δ�
��$�{�X� Yˊk
�"d>[��O	S2cևJ!�������b!o��j2Dq��/�dv����d~,���!��Ƞ�KL)�0֏���q� ��m��@�y,G䡃ldq:��s�[Q�6f)z32���D�Bp*�)�!�H��{��I��)��ԼMY�a@f�dR�L%e�
X�uo�X���T����1zN�,{��w���Hw�!���bG8v�~���ߘ�Aۣ'+Ĳ��:�ɧՅ�]4�}�Z��'��e�������R�7A��@�1�:�������8�BZ��;���%�/�N�HcB0��
p>�;��4����y
��U�8v����2茵��f2�c��?��e<������O�(�9��>S��+�_�����%+����.�&�!
})��R����K����v+`tc�9���%<x#C����`�\��^��5�Vz���8[Ÿ�b�[��N���ö�$����i��ۨ�M�A^��_�q�_q�5�Pq�q����Of�\W�X{��$A��ئSJ�bIu&_O����2��!��3	�$Zd�i� !{P0=A��疝�5���;욱�l�ZJ#�X��'���&q�3�U�
�ǰ�֐!w�w
��]�����
�&��9��Ò>��X��M���t3��tъ��A��Q��"�a�б�c&kѠce�I"��T	ʹ=Ն�zK���-�8)���~]�n�{�^�vI�����B;�6:"h��Ml�*�BHq���3G�"S|I�u��&B�#��8÷08{mM�S�T��r���0)i�_�]�� �$�<y
s����#�����a�u�V���$�E4|`�Y1�Ld�N~9^,٥��nuW���}�@ty,;[���b�Cd�ڴ�e���թ������/��>;e�e�}8:�"yk� 5T���f�4�t�vl��!9R�W/�@-�F��*��mFu_�ޚ��^Ѭ�^x|�A���+o��gׅjmp�1�ŋIj�9������Z��y��6���q4.�1gX<��e����@����Zi~;�%(L�]��U��A�񩺱�#��e.�nBqKI�š,�5��?�^���0=(NϩD���!���)?%ò�@qc��S��k��`�	Z��� ֬����_�s�˺�t8ӜK���C�=W�p?)��6[�u�j|B��	������e:��{(i��T�O��Z���~���c8 Q�e_��ܑ/�*!Xg�g�x���B�X�l���o�	�\HS�.`->�����^��FK	δ��J,p��Υ��{�w����hjR���:�5)��"��Y57���%���g$�ƙ��96��{E-l�2���Z|}/��߬�B3tl��I�P�����ƺ"C��%mX���¬�q[���F"b:(��(��+�-S_�by��W�|`��`���ˠ��D]xOh�y���zr�9���m���^k��oT�"1��5ٵ�mVq���W�d`x��%��YbO�}E�{1R���������;�A�v�	�j�W�,��� x|�{� B���:p!�aI�>�B�t`.��\�s̎�2���k�j�`n��ܪAW���T�-�C(���T�n.�.����w~T;�Y8�/�F�^Ș�ʉv��:h�;V�kʮ�}X1Iѳ�c��d�^H��%������v\Lo�u0,�����$N��,���o+VƤ]W��_ħ`��u�Z��m�a��ǖ5SdZ�Q�74Wc`ƵoЕ{KR	��y�s��!�i�qR�v�e$�Y��
�3���"�L���(�X�7QpF���ؿ���06{&���	�c^L�m�c5�U�n�?�w�+;�tp�w�z��/�Y����I���.�!�آЭ�H��Q)���+���,��ЯTx,>�/uUk�}|B��B�YUx��<�h�M�ꋀ�n_7��
<w:.��y$����X�@�K^�0B�T��C�$EGa��N�"2G��F.F�ZD�n�\�����uR�e�x�/��B!����U"�_��