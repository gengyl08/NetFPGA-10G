XlxV64EB    fa00    2540�bo8(2'��P�ֵԸX�b�K���֯�E�Ca�'�^�2��E?0G����@��9w\�g���u�����P�0��>��n�ųC���b��껹q��%>�b�7���� �0��duŵxZ6�\�u^S�
cϐ4Jde����X�H-��;g��S��hh:��`��B���½�A��(X���V>5�����Zz����F��f��D?<"Az�'D��gH�]��/�7;��2�����AK��`���(�z��*����'6�)�+ތ�;�q3�b:���/4y;[Z���\���mvnQ����&�dF������������T��lr�,)m��*���m<<3[�l��ҙ��O�P��B����� j/����̲��`:f��¢d���K��-Ep�q	�jpK�d[�YMT�J1y�w�S"��7�r������B�)��U���:�O������q<��V��q[��,�,������i�I͍������X0�^�~r��&��3Y��8w�Φ:^�9x_�>c��b�ܾ�$�����������s����$wX����U�P�a�*cd�n��Re�d�u������0x�"����>��Z�ԏz|:C�P��Х!X4A�N��/�S�py�����ƶO?���!԰aq��*��0�6|�"��sh�n�0ؕ��S��֚�u�ʘ1uY�'�Ԙqp\�~�|)ȝ8�Ѹ��Q3��˕�7fF�OU�s���}��u�~F��֏���V��,3x���Y�!��M�������**s4��Z��QzA��Η㈘2�Mb�YN� qB�`��P�I������܂�6Ob�ٶyt�a�Rz�-�Ū�&�s�eB���3��N� J�����9�1į�x�[&譕K����G���'!�6��`b��H�>5�P8�fꤼ޻���S���T���.p�/	���5��D��b����"������;-@�9�7� w��D(���9��~q���8i�+��� zK���*M��{��:����Qhn�~]q�/8Xw�5h�F/�ݢ
�WI��i�������$�����>�u�:�p����P�����`�g0����;����	ɈzpwX��Ĕ2.P�֢���)����N%�p���o�Q�e�b���xFݼ}�� �њ��3��bE���g+2ơ���Y޺��ݱ|Y�t�ػ��H!}�#���~�B��y���	ӲK����`2�$9�
�^��50�p]�F.�PDw]X�`��M%��j�U��E�[~j���Z �7���&�7�&6�Z�Yfs�"\�`^���)������&b���G�6-׏r�%��|vtv�rw�圊���Z=	)�{�I��28���/4ڀL�oX�g�λiڦ6RPS�xa�]e8cO��|��z^ԍ��D������̜"�%��w-!{(&�����}�w�D��'�{N�/R����r#%0�E�@ye�o�_uLk�\�N���ʿK�1�2W�&���I~f�I�z�wg�b
?ߎ���%6`�VG��R
��ҳH ��ECW^q�f�񓚤�7��22��L�w�p��_ڝ~������P�@Í��X�����$TIԩ9���8jd���'2C(�P��};XѺ��;Y�/���(�	�C�dhe{f�*C�	��8|�:n�*fe:��Ճ���k���#`˶�G������g��������~�r`S��Hr �l��iԓ$�l����x[�J���ijqrf�xm�m�~�O��36Ht�a'k�����v���s!y���]������?t(2ǰ|{|���L���M���s��s���mk/��_�v�(~��;�Per��w��V%2	�I��˒*��U�&n��+R�\�C��M�v�d������'�JE8���N�V뭑�ݾ�5��0�>��+��X�̀��C���4���@\ۗyٶǛX��fb�
���G첮�~��B"��.���I�f�E��#H@^�X�b/�0�r v��=�$�h5v�P�{�5�M��b�[��5e�[���B#1�9R#�3��{�4t���������|�	�;�O�80$�T���ɭ�>��nӮ�ü���.�  �N�x�	�S/,���ѓr~{&���y�����}�݊0/OE���h$j���������ﺢ0]k_W#R4�ܜgL]���S"�_�0:�/��N�������ġn�X�V\텔W3��	�����c�J�jm�)�Camr�+�_L�h�9Һ�䥆�W]%	��%�*��I���zb0��)2<I 5ތ|/���P��Ǩ�@O�)���~��V�W:7u����+'Y���?��{���^��n�k(7�_A��0�P���J�I��,\�\ 	J5��{��G��ϜJ�b��~<��u#gB��Ѷj�|7������{�+4$�^�3�ƳR��<^&>���� �� !C����k��a�05�Ӊ��Ӟ��8��ʕ���|�B�)Md��_(�e�]��l4��Eڪ����a��+W�2�>�Zf�{�d^�;7I�����.0�N��ЛNp0�2-���|��s�Y��OLX�p)��f�"){���:ә��%��T�/�g��w�?��u�Kh[+=�.{���[`s�\�c����fR]������f*f�5�Q�l�T����/a��<�RǛ@�#�S'7�v�Er��v� D��}\��g
С��,HXo��h�m#,ρ�_��	9*L[!C��i`5p�,�D�Vч
�W3�*�u@;�&���ɰ�5;ph�,��.�vP���}U�(qq�t�� *��lf�nB�����;5�ՠ�{����{З\ё�n��w�M6˵40"|�uzN�Z���Mx��Brh��x�`�OHX8�ؔ�5U�exc���Ė��ڶ�6g�2&���o؂$�몆��� Yi� 	u2C��C S�	4U�����$��2K�w�-2Ga�.9GHi�V^�Ŷ���iZ�����!�8{�)��L�{h�jJ+L/FBǭ��)|������s�~�q��NΝ��"���
@��fM�^�G	ҏ�Ā�VZ��4fO2ԕ@�)�C�b�r�̩�-��c��S�gM̠f�F�u,��toYaTG�8�[[x��w|�7�\5�<�F	���
��w���^H��$�kI/�D���NG�����g��I?E��Y��}�Dj��~˛V�^ �?a�9�H@�S�0t���ǧ��8�N���ݳpe��ʕP�,�	]#�K~�}jL[�t��X2}���J����[�\��h��"����*�>��ݵ�r�K_GP/�ov�E`���	+�h��:�V4�)�=O�E��]ʹ�R��au�����1�����\NkS\ػ��s�>��_�I��Ӻؗ�lb���v��!.I!���2Ÿ�W���r�R���ѵ,7���܈�%xfc��υkv~cq�x:�"7�(�BWb�z�+�A)Ͼ�Տƍ�xm�MM�ʂ�u��T>�෾C#	��nB*��>�j�֫")�T��9�����I�
�_d9G�Kl�1��9�"aI��u�1&��HZYj{Fp��/d�_8Jo�[�Rz�:X-qa��(� C����dm��q�k��ŃaBqS�a�{��Y���]/����V��`���B�g�!`m�i�����1.b9g}�n�#���}9�?T�f2-_F��P2%[�M�n�<�q���	�ű ʤ.���+���L�Xu�A'(j1��0�k�θ�8�obG��;�d�?X`�����?G%C��f,���D�w���m��=:	��bsxJ12��to�^���;~��{| ��� ^i���_Ƅ�SN�dND��ǅ����#�3��N���X�j޹<MP�����Xw��V�D�&��w�Gr?4>�g�f�S��-��n�/�;�'��Ƞ �ҢLu98AN+%�{��j��T��e=a������kP۟�࿹�"fK�7�n��D�����؋O�uH
x�@�g��9��៤ń�y�	;�l���̄�rI���$9��N��o�LID���2�Md�`�;��΂1��˾�; �g�.i� 3��c9���'�ޚ�=yL�6]R��\��;����OhZ�QO*�r�Β�'�æ��R���w�s"�Q������ �SJ�y-��3�#��r�k�&�Ɍ�����Ȳb"Ȭ�q��Q��Q�?�I|+�y?:59�V=+�����}�~��7�º�z��)/�g��ǸG[�s���<ygQķ]��-�1�;-o����+Z���_�gm��ڦ�Y��	�ȥ������s�yȇп�1�G�����R�M�
��+~����/����T-�6�o��������ȗ��au��eR~�u9,�2ҩ�\M��R0��\C�C��h��b��l(+H ��qx�;30���6�r"U\Ӛ�%!�b=b�?��=�p�r_��J��v�P�)��箵R�]���F�N{F���i���b��15�d$q�W~��MU��hY,ϔ�)�@��os2��8K�=,u��)�+#��y���y�ȇId�b���f�;5�S�c�F��(�OK���1P�<�EW/Ϳ����v��#!k�}����_�"OϩD��ul����Q��R�Z1C�SW1���3���F����<��Ot��hHѯ��S�j��?K1>���24��#,i�D�R	y���_�80���1�s��J�]bu*�K�4�����:s$�\��J�yF*n��T(�����vom�����H�.�(t� &��d<]I�u�]�s5ː9���Ae6�M\D.{'�i��ʆ;���<�^L*�R�%��'qP�z�4��D$ض��c�n��%���HoY_�D�A�`�)*�=�M;vFG��c׎oٰ�k1K8�^j��Q!�7s�pvZ�l�?�XP	�i)�F�8ř����^+�퀇u竟���ys��h���{��^��)ߗ��bw�)��ф��v�E�{	�T���v�.����D���W������N�*q�}^�v�_-���U��M,��2Ό��M��l���\YQVw,������a+]@���"s������e�S��]�@���HMY4*&݊�F����"�M�Cf�O�C�@f&�ޮT�r��s��
������� b�A*C�Y�"	��?�RL��Zs_�Ű+剱aV�ׇm�0>d�� %e�X�oA7*~�C���E����� %g�k��}���wT�G΄ ���w=����h����a.�����ycoω�;]�@%sÀ	� �`���1��k����D�`�`3�������튻!l��Hl���e�j:u��Ct�&Y��,�<����Q-�~�`�� "�˚�%H�8}����6u�;�;ަ��U���Yw4,��L��xW��E�w$���v��y΢�@-K��Eӱ�r����1�{	)�2oh��s����Hx��p�S�"�u�Հ�m�~��_@n�_���0�ʫ�w�$kTp��ޖWXN�Dj�%����K��dlHR���R���Q��l�қ��<{��[ *�g"$��{�'�^���\�ϦP�d���k۶�`�}���dr��*��XR��g���]#����$�q�n�}Ż5'sUi}(u�u���0�hbѻ۰�8k��&+�K��ݠ�履�_PH���������@�o���A����.��I<IF���'`��,�T���e����FQt�T��;I^���3���K�� �.���/IX'��ͤ����F�[ ���>�	���Aɟ�yl�󶠝�-�W%�\�t��ɮ{��˨��p�Y��2gys���P)4��� �)�:�_������;�~�4���_G�v�E�S���g#���√}4[��hl���z�IN�	Kz���b�i��u�Q疐Q��n�^2�8DϘ�}���w�(Ed<w>�pMI�f�C���ϦK����\��$�g5�O��)�p0�I�Rl�CөѺ?��g��K�ŜzbY�_e�m�!�6N�>�C��+��掆��7
��9��߷ب�ߧ���^��4�l��'V?��@�Q�^�Ĥ��:ٕ��.)u����B���]<��=��Ώx���@g���$�1��k�-C�"z:w6{^@��:TdEm��2ש��κ�	�ĺ]��5)�VF���)��_~D��r$;��,p7V��(����ց�S��"k�3���l+*O�3���>�4�������u����R%�Mi!/���S�f,��"KmV+3Si��PEPոp�����#3jҝ{k�J��Q���˓@s�m��¯("��c̵b+���a�;J�6^��?wx���LVu_�⛉�,V���?G��by�d�o������*X���I$1��Y� J�Iϋ��c�}�4t8���mo$$x#��ʶ����U����*K��S�@Q��٘���\�o�SHct�Y�p5w׌<��eډ�z�N�ʌ�KE0ˉ%�xR�D_K#�s���U�,�ٻ��Z5��*�� $��(�|#k��'1({k<b�y�=a�!�'�ñ�ܹM 26}u�T)i�J���vv[��B&$B*H������z�����y�	�Ҳ���鸴��3�|�W����>Z�K���TXB�C���rk˕x%Ԓ�0V������Ȟ��]�]c%�0x*ɠH�%��I�y���;c��9᧵|����9�ǣ�@:u�D�m�M����/J��=��C�+Q��c|�����,�MI�5����AGx�L���uQ @9�u�@���I�=;Km��֧�q�~D������t����GW��9���}�gf��;e$W��ٺ>�0-h4�8��ǿ�����a�|�&�B��!�ω;��2SfZ$�����!?�K�j�e���V�����O�^������ц�QYH�i�j(�^�~Y�hNa\v��Rv��_o�n�8�?*x��w}Ҟ��`d=���%5����P�E�[��%�@�t����][��jV�:L�o���W#=f]�N�FKػ�M�W�e��F�ɂ�?^3�^dŮ�'�02.�gGp��w��c0Se��}�#���F��&��W'뭰V��1ꩃ3FR/�M����%�i ُ�o�Y�����Y����m����V$QD�|�ڝ�CE?�	���.�1� �I�����ޮ?a�>&W��g?�����g%��RY��K6�M��\�ꃾI�O'd2N"��s��Iؓp[ޟw��1�C��c/���oY�e� ��Á�2~o(�a6	�K�}o�GO�����Q
�y�� /|�0��Z\�{S#j�FGN�
!GǪA*��m%E�L�wJ�Ϯƚi#�39�"qy��-c��������M�@}�>v�/W�M��7Z����O��O�Aw�Kۼ�D��ּ�fXU:)=�2)����ߤ.?�3�P�·���72�X�v	��vK˧�M�d��B/_�7���.��Q`1��9O�"F����,/ �T4َDب�p{,dA}���)Эeݩ�u�J>5���|�wkz@O�����u}��;����<+e�2���0�dih4꿍:3���ӈs�b�;��^A�91DO��-Gk�@~pk�{G��__�$��k(�ݲ��0���D|��\O�nX����k�.y<+��̃�n�����#e��ZtX�([h�@��O�JK�/�� QKH�
�.p�Ⱦ���O
Y��HMP�Tơ�`PPNڲ�v
�D�r�c�9
��k���dP�oaZz�r)_. ����oѢ狪�O��*Mܿg�_0�{.�m���u����1nRs�B?�����}�f�m���'�1p�8O��-y��A/:�;V�����|�g�3.���E�� Z�X�}�h൯*�7 K)�T�eA_v{}���+��8�&=��"PV�_Tym�*D���w;Ɏ�̱�7H�0^t�ǟs1G�m�|���q~-#F���M��ֿ��n[Dr2�K���d�$j�]��~Q�r��"z~:�cz~W7B���5F�t
y����K�cul�ֹ9A��{B������=ɧ�����2T����O����Q��>��6�G��ŧ#�L�9���cB 6�ٹoq�QEN���xPG'r�h��q��7����*6�� �?\x�θXH���z�1��Eʩ���9|�(#EQi���ĝ؋�;DK�a�v��K]�~W��Hz矚���k�F�/��s��7&���j1n,��@[�c�H��<0�y�J��Z��Q��\P{xu~�D���ʩ~���4bD�7%�/��8�_�&��oM=�2K�vȦ�@�z���*���4�|�N��d��[�䱗��%z�Q�K��4X[kk�؇_Zm���_� df����H@��y�l�/"��j�W"�����y���S�O?��Ӛ~e��?U5�uI (2��U��!�-1�<N�uޡ1��Ӂ�F _��sd��YЋ9D�1#���Zo��|#9ע��ǵ�C��'�����	j=P.6!֪�t�Ea�b�`�I�)��g�\K���瑝1G2�"ɽ�N����G��o
c�)8�<�����
FP��!�9BpKe{4�R�%&�iI,8{�/��(�X~8{{�<�Y����}|�k����4��*N�>j>6,����5��LZ#Ղ��3T�=���g���8��nj�6�G}{��9$@��a<[;�<L���hNj���t��4AJ9�u�M�앦��]�@UM��y�I3n��X�)$�(KC[h��2�$\;�g-�A=%8r�ss�V��ƕ#�����3N8KBIG�kvn����#�"=�[[m�\6�3��Z=�ލE%�t�Nw�1�Ơ��;
� �M|W���5�T\Sg��E�E����7�-����_��0ʬKɶ��S�c�hNX0�����ưr6��A��uZ����k�W�Z��sa�"��ީ��[�v5$_���i�� ��֖��9݁P+/��z�ҺW:��v(jV��O�W� %Ԛb��>�
"�Q�ɏW�fv!�}� c\���x�QA��M6��]��lʖ�K�����SP^��C/��v&��M�薳Q�Zy�؛����1,���������>|�A��|�:O�ⲫJ���h��8[G=�r��MA0�A��_h$���4�$U=�O�L0��[�����(�d��kmN�����t����&˃.8q�L�"�Mg��3�r��j
垐�U�=J1�XlxV64EB    fa00    2640�96R�>.A�JB���ډ��.�IyTN*/hFo���i�lw�|���<5tBTXWO÷-��3���`��f��)���Q�
��}u�^h���в���<�]�w�U\ۻb�j��>��QZ���r�iv��m
��=�!�Oa��`K�eL�G��ڻ��`�z/���CKH��l2���ٽL;���;�7��?�wM�6h`�bh�P�Hc��=�LE�Ӧ>嘭l�� �X��d�;z;e��x�3l�B ע��l������VLG�V���V�B�&���{���G�Ft����D$�V|�V��d-���;����s�,j<�U��Y��,�wY=q��X�(��0P�2eUŢ����Tq�cO���O�)�1f��N|C�N �C�/���Z��WN�[$vƦ��̹(I�����s�������ܘ�������zG�.���Nu��!��LM�R�K05�Φ�#5��u�h��O��AQ�z�<��v\��(�	.ZF�h��cQ����G��>�qF� ���s.������e'��T����ꊼ�O����cp%�_�����M�$�b$��~p�D����1چ,�s0���R�|3{�֗~�H�,LT�O�7���)x#U9�K�wc��gJ�x�m�4T�
�.U��g<�?�!�p�wż�Ϋ�a�����+�S~��rs-�q���:�Y�{TCy����r9�e�ub��$H�?��A'v�ў��_���9��ɇ�� qd�Q潴�]4�H�J����b�0����r�^�j��ޞ�U�i�����hԉ�#Hî`��1���Zǔ�I޻;-D�`��rd��n����~��%,��_ԅP�󙓙Hѯyv]Q����@޻��E5g�B#�!XQ�HG���\W��'�O����eH���'��#	�k���'!�4A��X�������'��'k����n{|���vY���?�%c��<U��K��v������F1�'y������dX����~���A�_%�����S�'(�":O%m����L�!�>R�����2�Ӡ���BaҦ�f<ߛKM��7�4R>Ew=��W��D_�Լ�j ��	N�%��Z��j��y,8�|4���
�ԕ�e��mO(H�v�X0g1/F�Mʷr"�T'm�F5i���e7Zo#�o'A��H�V����C�	^@�|�>eq�^�"�4�I���EhM�Th?�M�򚛥�"�$������b��o,�X�EƱ��/Ӽv�iV�#gey?��6d�a�hY����0EC��l�c�M���8�~��8h&-7�a=����%فo�����?�����T	�eB��i�i9T�#'a�v�~�}�(�j$�|�m�#�mW�7���}�Mt�K"@���˖7F+)�����-�d���ߓ�q8�oM�7"�_��NX�wI{�a+���Ղ�� ���� ��v�35�M.��O�as{e�s������	��������ge��#�Ćj������_D_q�"'���|y|��~0
� �Eg��}� @T�!��[�(���U��Tc���������k֜��S������2Yvɥh�48�jC��2%0Pm	�<���t����h�IRFEw�56J�+�{��$(ˁT=���<��M��͙d�[���6U�����E���e�/|}`�wQ3�%엫Ŗ̩��_�#%*ne��*2�	��ye��_t��L=�Iϙ�m~���2���.SnQ�k�ڟY�sy�����
��$��\���W�����1����G���>M]i����^���f�$��D�lzh��-S���&[����ܛ��$��+q�)8�����j�0E��jU�!C�:H��	[�R4�Nf}iƛ3���L�?������ē�Ը�9'���[!���O�0���'�'��h�x�7������y�j��v��$Bj�JhO���kn}zm.ۡP�l䬦���'N����"$��|�5S�l�}���>&����7/N|�o�f���K�%V�˝�Mn �ǚ[˯�$�8R[!��[��֧%�8m�նYK��ejjx�v��koMn�_��+�u@T寧����\��.H��x~���2��a��6p3�B����)��5�T(#p�'v�#q�g�'��,33���{eY@͏#�A���R�1�i����Z��v�P�ԥh�rX��芤YC�h�	fώ��`�� �5&�Gp��T^5S��uNon����Cq�pKN���#�D�|yqw������~H����)�,�+��'���sS5�=�.�m���`-��a)��:~�5h|�~���@<��N*RJ5T���T$7��A�S6�#�(��u�xҧ�I,�O�V-Z�F�ay|.u&��"��Nz��p��FY��I�4�d�������7F�����م�AkN���|0�v���
R�b�\�w�Fs6�[]ž�}�>9>oFO,��%���=���M�M�'�^Z�J��i-��Y^M������gP�5; �d�Χ�z?��~��z�ྰ`��������|z妈AHݽ,4T잡�s���ڳ�O"` �6���S�8�w�J��U�d�o�q���S��E��[Y8/Dh"�q�蒃�ƹ�rP���r��tMu�#��pn9Tt"o�����&XӢ�Buq�Ǧ���D���v��D�fDSk���<	&=lG$O�纩;�W�	{��o.�ȕ+�҈�]#�ݻ���bg�ڹ���[���@�9�M�ꬥcw{ydk'"�F ,"ϐ!խ�q�-��W�)�i����O$�Ә$Ubt��4���?��}��8z�K���-Kfyx�"o52�d�_`�8��Z)
"Gr��å�'�]T�D�NACs�S�6� +��!�)F�I2s�*���Z�'�3B�	��@Pk#㯋.���& 8;�]c߂8��02�N�u��n�1���{���u��a��P���P/��2�&�=�;Dv��������ՎdI�ģ�mNa%���,���SF�zj�ы�~Y��a.T%�ߒ�G(��q5�	(D	�z�xL#�Qo��.7���q����#y�Ï�+V(�����;�6����:)�U Y	C�ECݖ�&N't�R�5*��'@�8&�4.��"<�e��+�V&��+�����W��3+���Bg���h�;t������.
����Ėǈ˺n9��x�o�iIA�ƴLj���C��?�����V�c[H��({��e��9y�����o3��E1L��`���wj�'�a�im^���z�_��/\f���Mm��c�ʵki�+�j;1+�W�����R���Bf��QEM���f��P{D�w������drʭ�XP��nگ�6�9���:�4��J.7�$���	 �(.�ތ���DN^�f����?��{�l

Yq��W��n'�M9�"T�qp�鈇��Ҩ�n���i�R4��3'�����"��U����������&��+��.Y8�MSO���8�S�ϟ�s"3QR,����2b�7��dq#9�~&���z�iq^:�?�~���\��_����y́d�0� ��.���`M�cg�>�q�(�nտ�u')fH�"i/��l ���ս�q��uNj���~&� ͨu���0��.�$��iN�Y���W@R���>}����m��o�d��Q��>�����~ƘT��C�R��\�+�/�
o	�U����8MM�f���-�x�$����a6��yRY#B���	�v�Z���U�ɂ|.�4[��2�իUg@��g`��:?� � �;V�p��b�K� �e���3V��y,�F�o�fUƇ�%(�B���v�9���ލ�xR�E�Q{����ټ�&�h���޺�-~����w�и�vh�$DqkY�rx���'Y���~�z�(7�J�{���孉e���a#!�~�bq��$�~�}=7b�$�]����&�fHR�%]Fd<�Z��J.�����o$�5����3�0t&��{�ڃC����f�Ѕ-�ʞ��ے��z��f�oH��qx�W����O�U.�2hM�-��J�Fޡ�4��v��r&$�E2����	�x��
PV��1���D�������W���?56̩6�@m�W�@�vάI����	L΅R�&��ƇF0.�0�N���C�G!�?�MIR�y.���nOI;�vx���N�ی$�E����R�~+���_���l����m�s��P���p�-�VNWᵌv�����cچ@��aD�qE�o,�5��YS�'��í C��8K	�5�̴_�W���z�J�϶�!����r�:�`_ѭX9�� q6��lZ�@[ ���[�21&��N|�m����TqXW��D��gaJ'~r���N��PM��L��+�v4��O<S�z�����`�Wuc�p�%�����˹�>\WQ�l��x����8��+~�F���bJb��L0�T����}f�
�{@�[L�E��G��@2D=čh,�P��޳*����D�$;x�����.����u��a�M&�#+*�/I8e��96���!�aN*��dC�~����Q����f>?�;��cS@z��
3����QGb2��&�"A�+}W����|_��4�:��=�K��tj����������GM���`
aX��r�zQR&��F�,.�c(00�oW��7)#ps���T��FD0�3���ƀ�r�e��܍�`�Ë1[������2��%��5��2�DIS���R{�/=���Z��Q+��rV*2d���X�]��-��yJ�Q��SZ�����F$L�=-T�7@$Mސ���GRΫ͊z<���X3��� maK�S�.��#F���^	ٴ3�[u�jS�a��n��Ŀ�<��rŊ
?g���ѡ>�c�����ua�I��GR�)/��5�ƙ(�=a�G�{4�7ہ���#0�8��P=��L��% �lY-O�j���yw���k/�TnZ�@�A�~�L~?�ջ�b}{���.Z^��P�6y��P�`��0���TbٺZ���un��њX�Dj�L�x�{�=�-.Y�WdX�����+��,V�I��,_���ި�o�b��z�\�>��C�:9��O*��Әw�/��a�3�.#��Z�x�������Ya�+�����1���j�۔���-�JF	�O Y�o4��O�V�,�`C�#W��RPZ%�$O<��#�;���������7������U�6觋�2Ák���}��p��֦%sT�G��>��_�&]k��z�V�Sh�Qoy[J'.2w��/B���QI5&�aJ�b]��Q4p�.��IC�ZX��z��n!��d�O��Zf�1E;��髑R2�}�_j@�T��+G:<�r2��v,i�a8t���n��ݢg��o�����͓�k~T���ΨG�{�T��AH�A�͵��㖡*ȱ"��0�N����<���aZ���%nFK"-Z�����xZ�m�F\mS#ig�f�(����f'�D�?H���y��0(dR�v�����]�IfgT��PN�.�~`�b<1H��90<wy�&J�`qq�R��C�}��3ۏ+�8p��"�%�f�5U��M�� G�`"cF��Q1�3բr��̽4/=#����*�$@bd��o� �),X�p���k�gB��̾��{/��!�����p�Bd_L⌿�w��v�:��� z$��߳u ��z%[���;gR'�ˤ�H�p�$��Z�殥�uq-�E&��;�K�5@)�@'^���)2����74��Mu =3���cf�ǽ��]$�MX�
O<�܈�[������(����U,L�go|�y��>C񊮢�6qՖ.Z2�0�6Ԉa1 ��+^wA�c9d�n����{*��:��ڨѦ�g:J����58�� г��u�D#c��S����)bl����ϱb��ƞ�h�	5  h����w��ҫ�]1`8���\Vz�ϱ��d��������_�%�r.F�k����SE��#�	T�g.�X1|����Ԟ�<yOA��Z�����|��7���� �g���(�g��pq&@}�\� ��$]�\��<Q�*���t�{��^���IQ�:�k���&?�2/$ӻjkpg�=^���=��@��,��>E�<�����{�U�컮��(��W(,f�׆L�2���C�)���v��6�ҁ��r�͋)(����8A�K?�B��{��ӿe ��G��p@y�e��:[xB�>�s����]��̿�(4���M�{0-�Z�:�zs@�6�L.1Ţ��m���/�o0k5�t����!{/�����'ë�X�m+(�T�&�/�<�Q��l�v��M�@9�Z��ur	X��~\�M��kU)��x(g�����0��'?�ň1����%?����{�e��pt{�5�Y��^�|�����]�:��(NA�OA�C_%�ˑ_���oTx�ͥݙ��iwf��@ D���T������=W�~n�Jx��S
�&� 0�p��Gwqq&#���J~���Lo�_<����#Ew�:hO��͸|�*��}h�����X��X�z�b2]h�����g܅��:�m� ;͖xl����A�����?Tx��~��H�p��M�8Y�B��H������"��V����k>J�ex^��93զXΉ� 

沂�GW�.�= Б�� �L'�6l�@<j}k�!+ ����"2j����ޝo�%�%i��1��~�w�[�"�1ɺ�a�D����	=�<���^�<ú6�7�֬�h�;��;�3����Ei�oA�{e�
�F]Ou ��1�XwӜg�'ߤ�J�/�e&6�	g�|s�,.���hԅCQ4�؄�u��֬2�9���v#;�At�{������W��z�L�&��S���	����.�^�Ox�F��M9�I0Z��u/0�eP|'�~��qz��P��9\���]�~�t��"������9$�yU�U����H���
f�����z����}�$�Z��ƶn�'eBP�n��%V���~E+��c`�}���^���'����b9Y��Z�F��i��~W��@u1n�p��������N*۱���I�l�>��[�@ѧ�CNb��S�1Қ���+�g��B�{���͑4C�����g.�*>'���V�  ���`$ո��h��#<s��� ���a�g� ��Qɷu���^.gY	����qw����kۦ�fa�"[Z�~nI�C�i��1N,5l�{H��g�H\�/�QM�ʚ�I���0z�� �(x��[AS(���>R�ZM�z���m횧��jd6kv��{�O�Lߩ�~���_!��U<��jE�:����v����o!�A��?䆩 �n��7��k}i;i� �Ie��ftS2n�4#�𭾨���M>͌=���B���k��Ǎ*�Y��U�*1�B�\�N�S�����c�uLb֧��p�i�4&�X`b+P[p/?��"j�1�ܘ�}�C�������ۍ{�j1��( .����5Uɶ�꽓�������[��֜l��1�v��ʪ�*��&�BSM`G;�Q�+�E����ya�I��0f���
=KWѴ�!�֤aBQ{Wn�tF���� ]�r�
��'�A��h�e1�کz7s1�ބ��keN��0�ҁ�bٺ?J�&��aJ��u%n`��]?�S��������߉!��K9Jq�幊�~��Um��rE�m�!@��r&�*;uia����}� h�S�\�z�K�s�	�0Bz%Y�V���tK)���C�>�3���#s�(dF`8�����,��� �c���PK-���b�o�[~��!t�O�Z�[4eF��u�"�s-����o��Þ�f߼{�����LZ�D ꍓDęQX���t��A�%�Z���/�!���7��h�Ѳ%�V�3�x�>K����.b˖��,mUZ# ��m����H�� �����4v�!5��~JT�xO�+ӌ�~�x`���*��ҵ�b�{5�]P���]���W��;��b0��_6�+���|u��F�S�T�#�í�f��������v%�_�QS�CǮASuݹOM��4�ם;���'Dd��~�Ao}�9���+`c�f��w�5�ņ#�dK�C���/K����-z������N��l�I5��4$��ɖ�ά��F�XH��Wu�̾��(�B3D�/g��Z�����lZh���Q�sx}�҈���/�b?\�\y6�C��NY]T�I"�8��hu;�l���ʚ����r�G'��Q�b˚�+�����)Rf�5V�����վ�A3��J��� ����t����x�x�p5�">p%g�@�"h��Kݚ^kGjW_�z�"�؊��#�^L.7��Y)�����U�eʲM���x���(��Or�v������--kE�~���)�>N�|
w�����c�{h��`����=D���g�N���co�����]�:�W .�[t��`�?>�&�/�,���+��g?�6�C�~������xV\�t��'6K��v��;��VC������A|�zơ���o_k�.�O��%|pr{�͸�Tb��y���R��)���,��u+�r~�/{�����rV��9U,4�!W���ŶI�V�,"͖$Z%
���{2H#;25�	�1 g�)��v��w��b�I�v���B�UI�!��w��8y)�ЉԻ��\
���"-+(~5S�V�115��X0d�J��y�*cep�ps�^��]X�M�l"��K:��
�|��PZˡ��.�TO��B�x��#�X�n��ƌv
[=r{k〩�5���.�a��r/ -?��g�4�+�f��]���i�Śv����&9+�v,�� \���C��4)Ƈ��a�);��s 	���8�yh%��#cwY'�W J�I��Wc

��؞8�j�ƹe�zh��jF^����j�~��H+Hj,.i����qߧ�~̾wYy�>�z#�U����w�)��a���H�BBu��Y�:V�F��?J�QVج{?�.XF�U����r2a}�ۊ��պ��[MW��2�=�,w�����P�BSN�B a�E4A Mg]�'>;A��F��tF�7&;�������tT9�� ۅ\���pRqs�qE����2k]�)E ����#䌤�t)����=�Fp�����d����`�C��ɼu�:�6�]�H�0��>�ǿed��@J_����ʯ(2�3�dF8��Qt�*�*�a�hiO�j����EOOn��L���W翾�2Vk�Pʩ����L�o9���|_��-綷���Nc-��@W�L����6X[���wM��xA��FF�O��\��U�F�j���}�V���y�4�l�k�vʙ]�ݠ�V�{A/>�1U*tO���gƒ��Hpϵ��bH�'$���VB�}5Ts?���\[~��7�����\�S�so��Q��Y^�ZM?��l�T�me��m>I�F�/��%BF
%3�����K�����Z�6ڔ���k)�- ���JMny�Y����1D ���\�������e�@�;]l�C(p�AL��o����+�ڭ�16W�+f�-,��XlxV64EB    fa00    1fe0_w/�Z:��/�"\��%d����G��OL���f!�"aN��z��	��eGv�&�Rjъ�7��u��$+����*�:B����6���ހ�!ݕӴ�>t����r����d�ƾ�̞�z�(���i=Wi��A�� �2H|X�U_�>P�㹞�� �9����x�q��y����S��{�<�)ow+�|}�U��AW�|���os���<���0m�����R��yX�D^*�$�R������EXG5�(��fC�z���c��EX����F�RGu�Z�@�R��{�� �ܝ�fi�"�������bΥ\!I����B��E�9�Ļ�c��p���>V%�>�HC��.��I�៤�`8K�v�A�!ؔ
���&��n�TW��"����ͫ��{����q�Տ����մ�>���Ν?���Qj��.缷&92��Y�����p~tm�hS[� $�.K����Mt"b���a,�A����	��y<v����_iJ[�g>"�L>��mE�T��Nͦ@'9�R�]�D��:Gi���4MfH���_��@Ё����7��ְ{$ar\<2��s�mT�k�k�o�?�ǳf���B�i�z���@��!� *W��{�f��+�k&����Z[�� ����B�4�0�^$C�v*�xA:t	����2�A�ZMUS ��~��bً�Â�铳5��h~��`�����9��*1��/U6�JIFk��u>!��kj�J<���ۊ��^�8)W�0�/�UP) �E���5�2�0�b������/}l���0a�@��s´Խ���9s�u��� ����4Pn�M,�ύO]�V|�N���@-�7sf��=����kc�=�\���C�Y���QQi�?��� �J��Xs�l:g�TE�a����`�S���h�3��m�!�<���oO:Ud�>-p�eƂ��B�{wĄ�}9�ra��Ս�e�*+���䤿��W>��G_S�\��?r��I?-�*gp�`���b"��kמL�+�{�A�!O��㡡>4quɏ� :��H�Y��2- ���Y"7ӎvap-3�4;����Ť��*�F�p��h�0�ό�A��)!�.HT��,���L����:�:YE4�C������_���ΐ��<d�uo�簪�I��nn��
 ��UQu�o��`=WK��^��΂�2����ߎ��?�k(�����5˖|��r�ȼ�ڃ��*�{�$,�#[��"q�8+T�YŽPt�
!��sjFR*�y�ș&=���H%e
����8o������D܋�������V��PE��0��K<@�h��\qK�2
h��ڻ][�:-�rC�@����\+u�k�IKص�����/( ��N��6�L�[x���҉����#�7�p �$F���3{B:eg�nP.��[�L�U�x�N��J,�SC�6ɖ��踠.�W�'�!;���r�pFn#dU�#���o>��$8�c^u��m)G�~�@�L?����`!��М�tP��>BС= �fK���S��H3�be�)Q�	|�yW�V�vE�\��&�S��d���~��i/V�D4�0��*π��dwYV~Ty,��J~n���@�^�����U���e&4HvU�~��B���A�x�Y� � {�mj��^Ș����d�	*�f����n��tM� .��O5QP�6�Z1�%�ZF�t5�TnP�7�H(���!Q(��[��v�bI�1d!�P<5~�@��q	��fb���qW'}�oW/QdXuy4{WGg���\�n�0��j��� ��F�Dݏ���2Ď��e������ߘ/��my�c��ގ�����Z�ur<���_+J+E���Oz.� ��-�\�o|��ۥ��� �ˌ=<�)��zՐ���0��r�A���I������C��n��hb��J�e�'zdҔ�k�r�!
�s���퐿�=l̴,1��W^�	�;(��WP�\��_1�n�N��2�di��y�I	?k��[7���0���י�n f���M����*˿
�A�;��Z$G⿗��x�PY�-��\QBio�IxvK/��r�E��]�r�C�儎@�������喌"����P /J7�Ҧ�^�(��WV� ���aZ�K�[x�	�]-`'����ߓ�MO��Ɣi�_]&�Ε T�n��iw�r��ʺ�w�#̬�!�.�
"�}ȶ��w1L��f ɝ�e��f(B$��a�;%T�|>��6�u؜�K�t�*�(�<6"��K�����4_�|�� ��kb+�.}���X�\|<�+�{��<I��g7���jVE��-��f~���T\��`$���R!���;!��"�Ō]
��9D�M8��O@����x-N��A��S���'�/���[��#�L�B l{)mVF����*�pA�M��(���~-������{�:�Rڎ[�?�))���f�^Ho�����X�±DPH�S���]e��	o8�����g)�ma-RL>E�]�#Mץ�>���Vq��� �e�m"��`?�u� W�
�#IE]?�q���p;S�n�V�4�����j{�TT��A56�o���kj2d�h��<ҷ��3z��/�I��X�
n���kؖQr�Y^����&���w,���p����'���)|��W�����S�ձz�ݕ�'��L�J���Ot�� �q��v��f�b�¤���Nv��������� O�-�������h
�=���#뵅��.������:�4�f��5��?(�4�I���u���#3��8��[��`��Ĩ�����I��?��um]�Q���<��V�ف���H ���89����(޲Z
8��[w���^����hV��L�d��I$�N�J����֞���6ɶ����4DP���i�=Zl�\uR�J��l�|ʦ�O�o����4C�r��53�R�u%/�畮��:{�.$��{�����F��{��.�NI��#�5�z!QD��j�ͤ�X�'�ݒ��?(cSӏ&I?��N:���|e�����e��2~����ҚM��h�"*�T�Ovre��^�sO��$k[����Z�?G'�`[���<NC ��'jH���P`�l0��f09�W��G��R��~�y{B�j��6�➱P�}����斞�Q����E>ҕi�-�!�ϝx^��H��c "�9N�JX }�d�O�Ŭ�y��^��M#3X�}X~��̵�����QQ�����w��O�e2�����x�pFF������+�=^���4� .�t��Lb9ۻT�����zo�=2���� ���o62%(#��;Ʉn/� tiġ�O�d^ ��:��;��`�[�R��jx%�m�i��z��t���ki�����z�γ�����`��d>Q\�>%"y�	�o̮�ju ��0cE�q�D]瞃,�S�ܨ#���Qy��q~j���3](8�j�D��J2����oh.�2?��3/l�]d@���Q�h�޹�b\K��ἈHr�WU��;�AJ���W-���o
�����]���;�Nή�\V�.�(f5��C�{q�V�p��??�1 �5����5+�w�(t優��}8=@:�YP�<f�.�� �t$lmɻhl���S�����0�τb�@͜��ń>��3��r m|����~�����|Y?���³�s��z�"DM�����;R����$; �P��;O������MT=�s���q����"�D�����и@�^4>����vbѨ��K+�B�M�R���bW��ȍ��QxF�ŽX�k����,Y̑��  \��q��|:�%��V+���/��8u�v�����s@o��mƪf9�O�U0��~X�y���q��P,�[�V���Y
U��T=�τ�z���6��������,}��?������YJc6+�=㠠eF��nOk���= �"�w����?��5���L��� ����F�z�����&�k=�C}�U�8YU��
m[Yk���,$5J�w����x ��+�B#�Ψ���*(�IPs���P�<�4���_o�,hT(�Q��Q
��o�[h���D�8ђ�(xs�i_�؎�|M%�<��7�C,/�yM�
���6�9�ST�=oP�Ӝ��:���N�H��lN�����qLv�t�������ˏ���p��;JQ�D�o�Iܠ�09�}��ʭ�)1	=��/��Jw�1/�3��X�b
Wpd�`��]�F��l0;o�5�|(���Ɔ���R^�wĝ���1��׫��V�΄=��R�uL���g��e�鲭e��������s��̔�����Ĺ���Y �L+p��	X�$��`7�̴2h� ���D�~xH�@�ף�1H���;z��CyD���	Zw���Y��fq���$*�OA���9��mD�Z7�����bk z����s�{���Wg��V(������b�Z+x�n	� :�R��n�똊�2<D�Q�
���D��d1���L�äLJ�B�a]�0-p*[���H���56�3v[�F��Z�|�Ï��]���\;GUe\eר��L{ڹ�k�[�@�D���uww�R3I:�N��.X� ���M&y����4#Op ��5��Q*�r
/�U�8���m���!	� ?߂��^�]`AQ� ��(���C�c�����$Y��1���E�!�Sh��t�ΰrR���>�#��������K�<�iJ�ãw&5��8��D���
�3�->]��%���C��4ף�`���ϻ��반F��Z���f����Y�����Ha4�S��S(�e�Hh,��;�t���o]��TK[gč5D���dg:W��j7i�����KtY���,qa�Ǫ�G�&�����cBuص:(�3�hf !z����{᝱<AH�
UTP��M������f"UA�S�9lx��ݙ��v���
��^�{��Ȥ���P`�f���O��uc��Pm7��@�{A� )���:i;u��W��9{�L���A�F��[ىH�W�b~;���Ŝ��q��ڪ0��۫�{�,����~7ۚt�J.�G�S��-���B�#��nG��/��ح ��-�����^:6�h;8�;�T����R_E����/U�f[��|6�X�^�Dp*�r~'�����:��9!���O�FUNzn�!�W�UP�Q"������sK�f.Y���c��E�J�>>{����阣�Me��5���i��u��?��C�+��9/޵�'a�˧��̐�r�6'}֮
Γ�����u=|�z~��d"@���'��P}H�m����iR[Q�@��n��9 ~2�s���r�1m�|De �
��(�!mǇX���}��2["���T��j��MjG#t�޵�y!�����:jZ�E4+�,��V�\��0��^�+P�6�lȭB	G�ښ�[��>�4^�v"S�o��N�G�^��wB�0�p��;��������_R�M�Laͪ�.���ɻ`�q�@Xq�7�-[�[Ο�ON��g�&,jo�̒���y������s2.oJ2+������p�3e����l=)k;��$񝑏�Z�?[A�i��0^�a����N�5���	�ڶ ـ���'��E�H��L�U�[��J=�t�C=s�X�[��(:6�%Ӄ�ӛ�E�oƲ�!�K��k��e]����:��[I����A������١7t�ԧ�7q�L��k9�_No"��Nsi�s��0u;�C0N�޸��O���i#�[�s��t#�#-�wF���շ��Gü+Zj�r+�ol��Md�G� ��E��}%�M &f5����J+�U��#��ۈ: �w4�H��35b�#��x؊(i�UH�,7�A�1
��L���j��� T�ٚ��q� �O[g�1c���b�>.�|btߝG�=/��#e�T�6}��#�mq��j<`��ig�p��;�[t���Mu�A����_QxfR�[���9n;��[�>Ɔ�LAJ*�~s��G�%}���U^��!�*���;���(o�uZ� =��4�E�T�i�6 ��*���ݯ��l9\��-W��s�xLG>���vy��3N˄��F�rr#��Qj
%4{�0fE�`�,������#Ն�� �
lOR��YE�J1^��0S�e8/��4��Q�[�&���!#|��)d\'�jk��w�ST`���A[�7��������U��p:<T,9��N��a"�jಡť(e��Բ
'��?~o=������Jѹ.����5�K��$����|�l��bC�q���&�Cd��C{�<�%�k
~�GFvB_��v����t�GM�ث�S��_ʀ����~�N�� �WE�\�xB�aa�\A���/�H�i�|���)_�>w1`g�$ڹ�T�s�0������Gƚ��2�P��%}����_G������Apz�@����`
�Wo,!X�j2����>��z�G�zcks^����l������ G���oʢN�]�m���! x�*�I��^�b;e̛���7㣇����.��H�+��a+�?��y3W<[���ȁJO�N?��7�f'��������
��W�"I�¬�H5&�_Y�^#��o��杯�|�@�ʝ,�,�V���G�F6�� 	^�����-V,�@z��N�T�^!������[tu��q��c�%n*[���W��CL��K���W�3J��剭�2�M�ۢ���tc*�7-��Lt��V���e�Q��=.���]�����&~�^h�'����J||��wo�D�C��9��r�f%<h����_;&(�mߦeRS���+�l˺�S'�&&:���F���1o����_��,� �Ն�	K��e�'��П� �k�H��h-U����31�[��r2�I	@���S��/��ثDʡ>ɬ�ޱ|��/	?L�5!�I>�s�$5$�/d	�e �!�^�Oh�7i&�҉��l\u烟5h�(��R"��F����!{Ota���ˈ�_ Z�Cu7&Y��B��˅o}���/{��/vމQq��`�@�$
lqK����x����} ��Iķ���!���tw�D��I!�g�=9��x�r��]�VO|�\(+ú�<b��4����7��;֞��`J�p�nv��Kï]{��W_��#�U����?J�Y�+Dp�ձ�\��Hl(*��6�9�ab���y<���z�a�����#�]9�g<�g`�\����_6�9J��u�g��c�ⳕ ��H��HM�������RiSғN�m���^�(}�U��j�OLپ�Z|A�akE�ѫ?���q�7$�]0�V[��K��X�����Xq��kE��e�x؛+M�Nẗ́��X��Y�"�_�st���!��%f����������l� q[��&p4̈HU"������0R�V�����xB��5�?�~��VL�f?H�^���$�l�|i�SLͨ���'���U-Q�?���3�hx���F����W�h�e�J��r��y'�S}X��M)�հ�����k�d �o
!a��H�HK3G�r��$��2��v@�������~�LPoX�r	l�E�V6���Y�Qf��̑�"Tū��?�̪mW����*Q���Xr���e��l�9��o�����A	�*�6�0z���D`cD�ބ���8��j���ru���u�D��$\��n��$ïА`��u�H�=����R�:*�	#���u�x��^t��f�iZ�0ߟ��7Z�L�*�� )�"�݉t����j�AQW\�F�K#��Ԙ8 �}3�da^������� =��*����ok��Ho��݄(��+j���@sW�1��@<T|���X54|7�4��<z����e�)� F�萢��vaх�Y~�}N�[�w��}�b�V��"������O���Ͱ9p�
?��e(w4��̲�*iZJCXlxV64EB    fa00    2640@򴗱�K��]�r�Su��������k?0'əm��x��O��?9�kO�o{Ϻ�4v�G���Le��"Az��;�ڀ��W��B6�����ΒQ+C(�z7s���x�I�G��*��p`x�GX11bID��^��`��@R���,�=h#����lT��ț���r�kp>�]y��8�0_�Շ#��˷UJ��S�֫�x�I.k��/GB�J���������$����|�O�=�W���Z���5��[t� X=`dKYҧV-�~㏻�x�4M:.�"rr�oQe�����Ϡ�i��zn�4@,dia8`Ap�&글�-�E,��qj`{��Vw��ᣤ�u����U$�6n��1����Qm5�TZF�`�W��W����,j^�\p#9����o�/.�!^��|�� i��`">-���8W�73����Տj������0�����gy�~*}h�w�2F�.0��yc}!�x�/�M��l��������U)Ɓ��Md-�Vq����I��kee�Ďd�w���)�'�c�$��>d�;	F�O@,������������F�e'�q��;��Ӽ�L>�N�ڱ;Վ�R�Z��I��嗢n�X:dJ����6e��9�,Q7���Z;��Y�X�z7`|��3�'���t�����k@�c%���p7'���D��E�|��^�� �ţ�.�L�-�nϲ#!�J�{$=��2>o��Vr�L��a��E���'ys�`�_Ǹ��c�}�jƔ?�?v�������4�?�D�u�B)������.�� k: m��3�-r)�����&��&����#�L��N��I��f�[�Z^�w{%�*U
@�)�U�"Um��*��lo��B���q)��&���[��s�Hg��F	"���mfX�`�9��l�2$����a!
s2�=������n������u�H�W	��+�V;,D?k(��EP�Mf�u�n�bˈ��F��GS��K@��"�o7-��&fc�8� "G_~b嵆��7[��w�S˲4�����!���R�O=I�G.{X�x��/d�2�(�ng��ŗ���(%��B��0nR���A����0�G��e2����m�>�8;�f�@�t[��8W^;�ZH���.qv��9��0zw�:q�	�!����,.����sfOg[3Ȅ�B�I4����G��S���E�������ְ��{L�&"�%0�\�8|�hnp$Kz���� �y��A3c����;l���Z=����;�	���8 U��~'�g+`$
��
�7nԔPŻ!�mk�g�1���:a�}n8�5П~3V� �2�/��`\w���	����H,uڠ�9ņm
W��x[zOp�$���f��_�Y�ݱ��o����&�='q���z�����i�l��L�<�W�|m�z�%���
�b:Q�_'y�N� ��8V?��Ϣ_s���Jx����nT����9M����/�/�O�� ���"9J%h�;׏� 7�<̿V	(e}��^rYf�j(���4@[���sX<m�JO���l���Xm&��t�/ܨu-x7L� ~2Z5�N�~�휉 ���W�ƠS�:�o\m#�'��bA�s\-L�W��,C���s	w���k��̒���*V� �i��bnaG X�hሷC&;�}�{���n������YT���2ܡ)7e��i���+�<��Ť+B?�Z,�!�X��y/�˰@���{�3r�j�E������y;��mW�����Ѧ��1���%���n�*�+�@(���"����'����3��VRFL/0+�bKά�(>#cv��Z��,I}�ոL�u�1Vht<�;}����1�1�GD�~@N�Tm�b�� ��柔�\��y>���d^���<a����[�mMf�(+�LL����@׾�C�Xw(T:���F�ُ�(�0{E���)_�9�o?���)�E��eX?8[�\8�e��>ٰ8�ߧ�k�p,���z_:Ʊw�/�ƪ��bl�1=$���x��pB<Y��(���܈�J?��㡿�c�߭%~CY<���"���!����ɹ����؉�z���� T�k@�)%`\�i�i�h����
pt�/�7%�:]�ݫ��*}c����?I������	'�u5 ����>U�R��AS�\�c0H[��u�L�5���-@ƫKp�29�a6Y*�;��9 �i SF�q��Gx��Y�]� �"��/��5�G>2�
'LK�VR˼0X��%��)>�֘��!8V1ϵ�Z��B���I�~�.J��
����v}K�
FBQ�j��fN���tUk�SR�8�E���a~-v��R��]#�5��5�Ϩ;][�Ih�L����x�E+�5�3�\E!���ǳ<����(¶%��~~G�bD�,������I]���&s���N̯l�Y/���kV�K�3+�y�MhQ�$H?�sxfa\K���x�tU��*s�6��a�7�9	T`Fᰬ3��Ęwg�����8{�94�9g5	����E��
��G�1�}�Ty���^v�!�'�P��N�qZx�RG��nǉ�,��h�̖��z�ek_��:�!g)�����c���R\F�m��o�g����Iek���,�09�~��د�
�լ#��`j��K�з,}�]m*���`��������^f�ψ?},���J������_u��!_E"�聠k�d�g5	H<!�ʹzA�տGa�d3e�'X�9�)���Z��Td�څ�I�f�'Q^�"e��/��=���&7�e�˜r��Zc�+k�#�\�1�����pJ �:�(;A���l}����E����?��~���v/��~��X�'���`��%|e��X�f���R�屆�6vd���̿�V�0B��J9�C��=-��1M����v�Wj�A��%Vܣ�C��mՏ�x].t�W��*bk�胶�ҭl�<��s�%�RN��aWcgq�����џ`�q���=LuSx��$p+��CW��y�Tk�˱f2��S2���H��(*�Jr$��g��m���#�Ȅ9���`h]�o�_gB�(X�j��I#3/|s�gˀ�g�����<Ud-�/����EZU�J������: �Q��le�gx&TK�H($�V��Q�����Dk=�~�������K��b�fI}����<�wSM�SJ9������_A�\��E�v��#ja��B�#�q�V
��x ���c?��
�%�˭�ҍZ.R7`}!�pq�?��:���B��h��z������z��{8��Sv���ؓ��M��a��+[\�
�|�y��v���u{��p�IV2�Ąiq=]��.�=��֚39�2ҳ>�0��Ý{�A .s{4L���k�?E�P�s��<qK���ȎF��g)�=��<p�.e~��<\g@b=�m^ �i!���oIŉl��=t�TREl�8]�Y�%��h����� c�\y���ǭ���\~Im���W2~���� ���r&���]ȧl�l�:}Ğ�ӊ����}a<�@�=$ۿ�vZ�q>��'05F���^b��R_!�fs�6��Y��t��z�Ci[;�4���	[�:���!�}ȍ � ��k2_�]�Ö���dT�|�\S��WTN���z�%���׎���~��֦�>�`�Bƅ6{�������XNh����
��r�/�uN��,ˑR��m���T�Twp���Ir����4/�n�T_�!�j��ay�匙��@=� R����iҲF�(�~��R{]A;>4�!d�ۚ¡��K]�m����̀�A��jҝm��UB{�#(��^b��t�d���M�IG�_�ʗc��j>�?G7(�C	��� b	�q��8NJbB��3��Q�2U��tr���Y
�x�ow���<�EǬ�*c��Xe>(��bX�Y�U�<}T��!z����se��~�p�2uf8tr,�1<��Rui\tjD��h�6k#l�`�S��@���u����K�HE����
�c
�N����� �g�g��`��Y3�	��g��m��,���
�RÚ�FR�Qo����O�����0���i����o"5�O����ܡ֚#F���
 �^U��~,Ky+d��"K���<�I���O΂�w2"ɬ�XqT,]\��!��Њs�5�(qC-N��o����AΖ�T�g}j@�ʰ쉺�H	�� !<��^��kӞ6F���yȹk:�:��}�7lz�6�Ʊ�A�`��}m�(�4�&zm�i���4��LŞBp�
cg�s�լ�	�^pN��b�^��aZ9Y���W*Su���J���~]wV�.[D�J�ጢ(V��u��:*�0��l�zU-R. ���?!�P$y�1(_��I:��O738V-�$���I�1��e>��̨P�zp�?Z��O����F�nfP���Xm�����2���8e�Lߥ��5)�G,f��-�V��/"Z�o�G66MB���Bd*E�>;Y�����2a�m]3p�I*�Ձ�Ry������T�NA����&�jF��^���Mf���TƏ��ó��pl�#��
D�N���F'����y+b�cKvN��_Lv���	��dv�w��ʡx��*Kj�;lyF:^�M������)@���onϿ���՞���ޢ��&������%��6�=�{��=�z�#�J�����ɹ�ˏ���l�z�@��C���=I��z>���@"׀.s9��z:�HܼZP�~;=��L�����k��W@þ����n��Q��i�:�<��5:������4�]����U��Օ�" -��]�:�7�r["ͳxdq�n��' z��YY�N���T݆>��w�F7,�~�6{����b�c�O��[���� �Xϗ@���_�,A3�
���?[+���GJ�%?�bH��h�E,GTʂm �vt�Hfy�?��o��c���Eoc��9&��cq �Jl�$�y�xg����y��P��AvJ��Զg)���O�>/'���c;\�D��쾠&�J5*��j-�5H��^ne/xN#���u�
!ٮ��o�_0=��ّBa��II��5�B��}�쥘*zCq.�I��'�C���.�q3Q�v�Cˡ�g����;5*5�ŉ�]e57�v�`��f�!�l�R���N;?�S��ڜ���#�FD4�O�ˠ1㡛����'l�.�-�?�ԧlQD
8=��Yk�x��^p������hD�1���`k��K�m���QC�x���T2�H���0��%�ťp�΢�9��kdE�b�)��|f�-��j=:�DRK��dx��8�ɗ9n"L����ϛ�uY��M��!�T�'U
^-c}���G@����M@|��Y�e�@�����w�k�dǂ�KԜ�2ҟt}����Dx��]5$�c�����q^t t�MWE6l�t�Iwbs���<���!~
��,`Q�byX����-�"�ۅ�� 4ݩ����6i=���(�aW����<��a�zn���,��Q�pM��ʩ�w��Z9�ʇ�V�"�|���y�°��=K����:˅K�����A�T	c��WE&$oN[�BW�5�(K`�n̓�T�4��PcM!O�ɒ�8Fqd}�Յ��å���#�ѭ���<�/_� �Ψ�Z���Ԁ�J 4)<��$6�9u"����]o��6H����μڽ�֖�፴両H�6��9�� x�t�z;�כ�J9�NM���C5R���h�c�AY�4#�q ��Q�p�>Zg:Ā!��V���% �q�U>�
��\�ލ�~>���L,'�-�p��TzF�ߴ�����жX���:`X�|��'sJ�(�0f�DE��ҫ�TbW�_79��d��U�A�_9���e(�+GZN�X*�.�����6�KʖT���=�i�
M�[|�^%(f� 8XV�3[5�jJ�$A�v��/����Xq�
�{G�4���蕘��dl^�\��$�܁	Л���-B6�!��&�ô��({��������^-#欸�=�r>0��t�TeC���$x�S2����@?�ݧ�(���-��j�6���:�`G� ��Pش�:�.��������~f��fe�`p{}���D*�����B�',�8p+֣:���;z��\S^�g�΍X���_3���T����yY�j���ذ.Ώu���^��6j��&�o�i-	"x���"��ϔ���|��)��
D#�yRp�XyM�?A:��2𕋓쇧Ȕ��]@�8u����CF���a[K4JCud�����T�;Q���N����j	�џF-��'��#V�>�����"�j�
A��211�B !>��k�o�v�rzr%e��r,V�`��vid0/?�[~:+~��-�n���Xd��͆uG�&��P)��$n��O�����45/�\j�|P$NI����Ȩ
�OTX@͵�k}@��+�:�e����ASIT}L�̓���CZ?n�a�'X�ĳ�d�{�`�Ɖ$�ܧ� ɘ�ڄֵ���`����"�xo
Ü��8*���Ѻ�9%5*��.�dnxV�im�r�n�^X�����KM�O#˩Z�*���R�T��/��m�!��@�4R�Rٞb�����D.��m ���=������|O�Tk�`���b'�����)�&��دgi �Kxn	�� �X�'��g�u���s��1NgD��!5;@���8n�F��qX��1���|�fZ��� �=��_��U��02ȝ��G'.�sCӓ��uZJxB�oo�-~7M�[�����4��WwRT�`	���̙�fb~Ni*a�.'��o�,�# S�k����@��均.o�����پP"�ބ���̅����;�k2�4���%������qov��1Ld����G�O:�m"� �<�\&���r0Wo�����1����`��쟄���E�D%����r~��� �	*>������'�M�uy�}s;��K��.��p� Dn�M#�gRފPSL�f4����*����?�o�w�ҁSObr���?V{�/k�}�����Q����;0>ON�Q�b��v��)g��0�v�$R�F-d�Z�x�ð��'�+�a$<��sw�
���5�<-��4��r�*�����L��������*��S�i�iWȰ��L�s�vc.|96�!�ꑄ��i�H�A�	`�/�yF�F��Y,l ��:C��a��gj�1\n�Π/Ϩ����Ņ������P �@��o*`ͅ; 1��k��UuØu��áHvY�_0��Z�TIA��>:�3���10��4��l+����.��-�`3��К$}���TS�q�7���ZX�j��g)�D�QQ@�C�e���7`lпYD9S��������T���T��Ҝa������2�G:���@��@�ln��#A�,` C�FTʧ�(̣0ӱO��zb�1vd��X�(}�PP��iKb����@�N�9�{��|���(~��!�6�n����t&�R�x��D�I�'k���L��C|�����h�z�f�$%�Ƒ�۸�p>�2B�q�������P����w:��qx]FAB�e,���KA���%��R����y���
_�beO0 ����U�ܥP���>J�S��<?�~��Z��ͮD5"�$��֋�'��]S�rC���a)Č��ܮ̏@(�J�o��`�&j�i���g8K�a����d�I�i O�K|#����$�iτ%��b�#Ŕ��f�S0��=��tऽ檋��d,!P�_G�A����%S����"�1�ﮑ'����e^�8`�?ɏTU<�0��?��%��Ⱥ�?��X�^R*�*[�	'"v�t�����։Ƨ錪����R�13�R���Yp����OVI�"��q씧�I��v:*������,<Q!��s�f�wB	Ѐ�n�p^��(e�%��&}c�6�CETQ��^�!d{ʯhf`��N|SI�t5v�ʧPm��ҵAG�Q���:�l)2��2�����Iy�ٵ�jOǉ[��%O�p��͞��'�Z�O����;���M�C6/���a�	��x�����$�7+U�����>ԓ�O9��*Dz-_L����z6�T���h�#�ɚ����A��+-hAc�������z�_2j�*ޏ�h'�����Q����څ��#�N����N矻M� {N�m۱�񱬿/:q2����`f����RKƸ�M��l����mpBr��;���"?�݉Ĉ�*��x&3cjػ_����ԯ�6��PV���57©y�_فr���}_��S�p!�)GIo�!��8�.[w>�,�6R"W�K,RX_��XX�ȭ����X���Ul�P��1/��o����0�ֲ%yD��,�~�����bT�.�W�JF�~�b&��/;c\wb*���	A[@�������n7�S��=�*�G�_�*�����?�|�S��^��b� \�[�O�sq0T��3�9�jz�5=��{s���)��ň�7�cOۑ����7�q��a��(�
�4ޅXw:�]��Pߗzϋ���D@���~KT����XM}�o�/���|UG�Ї�6H�t��uj$W����]����!G�������6)/$��� ���]D0�@��,H(g&ҽPy�	��^J���S.��=�/�ÿC�IXb�*8C������3Tm�Q�#k����$g}㡌��vD*+T���3���K�A:��vwG3XQ�M�}
�N]��m<-K���O(E��{Yx�:r��Nz�}M��C��RB�Uܾ��?�������6�_�UC�������6$sⅽ��-} �6�69�@�$dz�헚E�����#�F���%��H�̉RR����u7�D����C���74�R�og�[3��pJ���g��]8�N}�H#����I@�
���ٳ��ç�
)Osg�ԙ���{V�[]��x�B�M=qA
�|ziH�2�R�m���;��X,�Bɐ]"��� �
�htPWV=���@Ѽ��'n�7�&�gE�4�?k�:�pKP8��ِ�@-��?b�m�ʣ�"�r��z��j9��d��"�Ek�!W��sJ�% M�<2qќ����]�9�}��ڎ +�.� �,�6�@�k�F<�5��5��[���\�<$�P���7�MK����<�w��L���k�˖0xi'u�����^�&�7K�Ϥ�+J}���)����Y�9�����{Y�D��y�4�9Sκ�mv�*`�%��+���i+'�.���M
)d��K-.��s���V%��}��'�^�����|�u�)���B��~m��Ȳ0}���ݳy�5��No�%_�y</*ʓ���&c~г2���~��D��$�q?��u�6�)���*���YV���b�� w��(�D�a^��>ͩw�܉��qg���A\λA����C�[>)�L�>�l�h�Z��Hsr�w ��j�r�!�����E㳿��ӌ��m-x�:z��_$��Lxd�^)>��4G�:s=�����T��}�0�.�XD%��dp�#�S�/���>SGS3D��}���R�/�rҤ�e���c�<������״j�D�C�XlxV64EB    fa00    26a0�7��`���:����u���?�����՜�+�W���0���`��C Py�1Ds��p"�\�Q_zυ��Yn�T:ʰ��W� ���vX���\���j��ʸH8�����
�9��_`"��Zq`�p�u�P�Ţ�#��������C�
���/Ϣ�	��>-C�����%^���'j������(���� )��O�$�5p4�4�+Œ�~�nG�u7��;"ī��2{.`Τ�����Wy'�f!��܈�翥�# ��������HY�r��ڿ��� �X��9���A�}EC;����a�� �"
�|��9���҃�ߡ�	�Ӂ��.�d�"O�Ū⛪��pK�8��]���?���5Ug]���-].cE��R���<�8j�f�p��r��r�-���`����>� ��]ib|`B�@����~���e��
/_���tyå	����$���'���r��u)��>���6?dZ��ؤ5�8Zh��c4������K��J�����9�$�eCJ>����Dt闉��B6�#��:h8���\��_
����e�F�����r�6�B9W�S��Ih�Y�@����W��A��m�H���i	�� �-ukt�E�i�ю'�@ҋ���k��(C�]�,�p�ي�YW�C�N�6N���w"TVs�H�� ��J�$�/n��=\��'ם9�R�p����9��1��3�lpT�i�K�I����fR�)��0�o�?�S�հ�L�'g�c����4�̞S�؀+`�3��G5�a�:��?�� ��p�۽��sP�*g��R�[U��J�S]E��p�
����l-}q�vS9u�0�\Ȓ�C��P#6� ����|q�
(�$�O���s��Zu���"Dp����ʨri�4;��"��=w���>>=���/��)v�X?�ͨ��gPj#��.&���ī�*���?��O��ii��K�kY�Y�Å-�)��7����O�j���~���u��q?K1�C'�{&R�~i���J�}�9�O�lw6����H�ʾږM��t�����`��&��C���Z�ܪJ�a��q���kB����9���XJ̶�g�,�'c}�l�L����@�fR��?(�`b���*a�����CҖǏK�l�=T�|"n��m1P��iC���|S�|.�{�cI���8�;�0I�G��a@����ߡ�a����b�!i�c?�ǧN�5,�ۋFq�9��R""��~���0+}���wX�����RLE7������\_ꖄ~��m�A�m�kG*j^�q�����9L��>�6�},���#b�ガ�#,�ol���_���2E��s�1��)+�C[ߌ���uwqp%2�T��}}Fe�y�C
#����>��r/�ԫ���P��%�`�?�0']8������;#-�HO���0@���w;�#���g�r/��r책�/o H��(���g�z)0*���G/���Tg/��es>��ܕ��&%|D�3�7�	H�0d.�#��9��/m�Ay�z���D�AfQn-���ʡ���wt���$��@��N}�����$K�US�HX����������ɢ�֏$7�5ٍ�5=MUi�]���@?�8�L=b��i�$�&�rHw2VSF���w�y���)͐u�U��-:�\���n�VQ�h��衶̴����ĲN�8GF$��]9��v�bLd����^d>�Kn�M�1gCr��L��:�`�dta��Y^p4���.��~��4�,�~d�o����"���{?`Hf����E��G0T*�6avQB�{j{���0�W氐������95������^H�ut�=^`��@�<��Pgy�];�-Ҕf�>H�i�?I�ƷO(��*6���M���R���Ǽf[���3�
�;�]�\d_�7}**���>剝�)ז8����ݝqQ��
3{�	�vBE��q��~�e:���w�<u�;��y�Ur���wd	O���ri�#�=��}������K�ĺ"�����F�~�)b `��z���\,X���wϯ_���r��G{�i�rQbZ��4��dG`��qL�S	ݏ<�3���$ursb���,r£� py�y�7�K\�KK��\($�i�&u�</�7qe�CQ�����hF�T��s�g�LǙ�Nj�
N���}��5�NAD� ���vW��Q�@�j+��$�o�|�'�bc�����[A�m$G��K	6ۘC�{��< ���M`+��1WVy���@�D��Gj�sW(m���Gk�]���
R\�������yIb�SQ�fg=���Z���sO��dS��=	��㞪v��ݩ-�hf�0;j ���&_�v
`M�31pMc��56�2�	 �f��Tv۫.����&F�|�l0o�!{����ӥ��e21���=��V-��܄@#k�"�����"�- �*W�Z���[1,sMs���L�_��DX�
,��d��bT������9�.���W���zF�`Pb�D;(Ly'r+��T�֬��Bj�K����2���_����jQ���.+p�̹+� ���3��	B?�5A0W�}G4�Q�@�qb�7������8�6 =�π�~�	Ky�0�#B��N�e��G.�ԑ��U�= ɻ
�=� ��s:�u�6>ƫ�zg���j�:�A�e ��'ɸ���4�J��}�B�쎎�γt��Dk\i����Ǧ�ؒ��M�v���� �vӱ"��`:�>}N�
9z���p�6xI[�.�yٓ�vń�3)��&�1�z��)�C%��V��#�
y�ncU;� ��0�j�;z�I�,�̦xpu����a�*8���en���T�(�9��b�[�8�i+r�~Xv�\���0ν��ܘ"��F)��Z{хq����?��	���8�M��'�����p#+�*��y�dĂ-�D�?3[bZ�PQ�t�_��C������Yӣ�lg7��p�~��|]�Ǳ���ZI#X�������}�3�_X����W_.r����N�>_q^�R1�#|͘T����ܹ�hN�t�gˉ42B���2}ݨ�HMa�sv�6%�5�����m���80�~;���CBHY�o��G��-��lM�m_�.�jyrg�,�Нqr�[M��)��޺G�AUE�:��&cㇵ4���E��<۫w7��Y�f5��6�7�9T$�k�)���ZY�n5�oBtԦ�J�L�Hd�¡hJ�I��&x�rg|uw��\8K��2�7��i��1r���:��D,�#|�N��A�0x�H�D�#O�h��ȟ>&6v�au{�;��w/ޒBW�O��!FK2Q%p��ug-���U��;*�:�C(�a�c�u���I0`!K�Hxz��� �2i:�6~���0�+B]��?ۀ8�x��Uo_A�W
�VͿ+U̶�Kt�vWM��b�ō>�e=��U�I@:�wx�Xl��9m�������(��;��jJ`T����V�%f�[W�R%�˦Q�5�A6�:`����B��V�q�2_������b͞����"��(0�:N-*~ØO"'��=R�'V c��on��+Yp>/%�3qe.}z����7�����h{*/Hjl�L��7�EZ��՘#!��fU��y=+�_�����gL60YpֱA����lA�سT����fIuӨ����%����*�����w�KXG�e)��:����WSF��B��p�dd˞lLOk�X(�\}������O��H]d�}'K{��BS)6p�S�}��rx��A����<w4c�i�;H'��G*7smt������9p����S�8E���D�/� ߏ+�_�'��z���f���0��e�r�lk�w�q�MhX=�M�|H���mU�
�6��n�2,b�,Rr]��r5�\��Z#C`Y��%�H��i�i��v�Ei�)�qP���X��7���N��M��������"�OZn1Bd�6q���`��3��g��4$48���023dt�㘄Y�G%/>.�H�^(n��`-�k�r�v���P����x'~�b��ppwٱj״n���jj�3�����D�[�5H
TI�pI�3�?a��h/6� M:r]��q��r�S�~]98��KA�_����$�z~1Xk���ܬ�����iK��
 �V�Nv�a�/��2)�0�(��Pqw��r��E���I�}r:�����SS>��i�
���8�7�>�$�\����(Aɟ��ӂ�~�$�V��n�<�b"S\@��ߑ���2X��(�{2ǘ�X�G�~;���8���Dl�EI��_#�W'H����x��<%��w�D�#��Ǳt+iMC�&b��[�����rev��E�U7���J���bL���`5�'Д�p�6��*�7!�2�����������E�J�Hѷ�f^��	��к�F�\Dp#^}K�W�M���pE���9�1/ԁ!9�՚����U�����w�����@���GVj��|��AvO��Dx����.�C��z�S��A/;��UP�q�����<?L�Ia���K�ؔ	UX,�מ2��>L�/@c�l/�:�x��iU���K^�'ܱ��Pҙ5�Z��2� �¥�M���c�e<��$����q�}����X&���:E�]`�t�\Tٛ9���L�f�6���0�"�j}�l�p����OD$��{m��������9��K�`)���U:3��&/tf讼 �:舔-T���7�V�8�J#O[�Zd��w�Q��$]�	U���8�6�@m��Ø�g�
އ���XmH���~�1
S�)f�>Vޕ�N�L�4�\�.��&Zw�Ow�B�	vR�$ln"�o�s!��ۓ�n����8�+rk�3k�H��B<pFw�D"34x��&}��v�E��ل��TU�.L���'�{?�tv�L��)���+�0�����������?V�(�M�}aia�¬1Qߎeոfu�,I� �{���8�����A�z��`���B��O\���j���n?�;�f�5r�p@��Ǐ����߱7ňKuO�
��<��Nu���P��FF�$q!�W��c��L��M���H�6��O)�ق���ܩ���x��(>̚Pzt|�-N��=:˯���?�P�v���t*Uϔ}�;:tY��8��{|������1����t�ވ�H��dO�2�Q/.k�,�QµS���A��]�k�S�jE�<4����g丁��b(z�{f,�z�����>�K�����>��cȀb��h7^���M�j��=vP�]���\�B�4�q�p��"��`'�]�k0K��-�}+�N�'?A1�(\�rTt����;&^FV6^a%��Ia��d���'�˨�w�'?�4��<w݄�E-�<'�cI�d�򵿱�	�l�;�ry�K����X�?7�?$X^d�c�J$l�h9�69x!lW*#��lA,��Oΐu_�����;���m�>��(�<!vG�Kb�@t8�2��{t Wv�M�Q�q�^��9k>����`��>���8�|[Ц�ڊ�nrs=m�l��}Qp���z����Y���J�$[�vG+�	��x���ڂ�h��3_�<$UjWW��}[�l����m�hIԿT�q��e�[F�+��I�����~O��`�W&|8w�G�'43/3��a��c�	�	���������z_h�թ-76j(��{���n�s�oW�}@H���ӎ���P���� §/U2��
�G/�F:�ً��1뀊8�{/w[�#Tֆ�9��r7D��E9b/�Vq�Ĺn��C�%I�^QĞK���Px�Y_��Z�,O�Lc�_��c�!��<��X�׎%M�x���3������2��J,�Ī���i<D��v.�w��H�!�u����8�{I�V���7�Qo�;���+����C��1+�o�F�A���}�����.9uO�dw�5�U.om�-b3�n��[�.�j|�>j$��y��]�j�b�V�eQ�Yw�x��)�=� ՋO~���$��>����*V1]���h�oH�߈͋�k��SQ�Qf�[x �(!���1���Ҽ��������\�S
c���A�(R�0�� ��LU�x7*��V-���o�@9�D��.�~#�/Q�0��H��v#��_�:ٸ��Q(cR�G�w87�g ��*J��|�q�{�zI���q���&�H�Eo|�A��{~�(Wq��B�@��1L�ݴEqw(�!Hr�6�3!tIë�f�"t���L��\��fB���Y��ב��<%ѥ�ry�WUx!JY�a�Y�w�d2��F$_��p���󇚯��b�r�)1���=���n�9���6#��9��h���0����&*������\�-���n���oj��ys
P���&&������V��19�O�w`�������ɑg���8b�!���d8��:u�n8���=rܜv�!��)���ـ2�؈Q���[��@Aa�K���@��WiK��i�6SLY;�?9E:$��.=�J~�_eo��k=����:ܱ�j���HyD�i����z���h����ą�4w�]�! ;���T�͎����{�ǡ�zE��e��P����q���`��No>�o§h��!��JaEf P~�r��գF��bY6ΖrOc��۱"	V�ܢ����k}}��ǠP,��i��_��.?�j�%<eחx���z7$#��X������؂�?돎� cdV���?�χ���	<;j��J8����7=j.z�U,���r�.�Xp��*znUX�VD'�Lq0�"��]��Ո7�r�:��훟7i9A��VI[H2�9��o��?��8۩��
|X�Etw�/���0u��$��#9��~�4����ǎ�Y����:�5��Sj!J��#n�����sݕ�vH��n�p?t-��#�|�j�Q��)��iRC�����\�(#�r�,��2$k(���j����޲'��p�-����X,3P���ppU����Y�d,~�S��El?(�}ր�� �����-�wb&��"�|e�i����n�(g^|�:Ϛ�2�%���T1�EH����m�f����]�t�X��M��S���YɆ$�ƕEFs��#�Ȇ̙'k�jx�}ڝ�0�H�l%��/���|p�b���Hn�7W,�`�\�%n���؂O��N1P��4�(��	Gf(�nb�u��x�`<�
0���&9á�%�l���nU��Gz��Y}C��Jz?y^(��� .J��a����3F�?�;Bā�SH���!gY"0����}�v����Y3��M�H�,��$�½�R���.��e���-vS�����YW�I��D�S�oK�QL�B��q��m���Ԑg-����6��1������(	�.�<�_�C%-k^|�*��}|[��=p���O�A��ԅ�`$\"Ǧ.�*�4/rͫ��=�3�3#��G�gnßx�kJ��%_ک�ʑ)jL��4�ChE'��]��T��߉hsa-�r_��������Լ��-~n^���3����|Q�����v�Cf'�?���w_3n&wY���G
��H�Z�3b��-P��������,�);A�\G�B��w��G!XfɬT��i�yNu���,e�;c��z����_���
�o��㥨�V���&����a7�'���D4��<�W���Z��\\��V�͓��E��)^�R��kuݙʓ�A�@��V�jGO��FᎹ���TjT�"��+/��JF�C�>�;#FX;�Rn�)D��)G��xZ�N�nq�E� �[<�^��=�1��95���_�j׌0䅏M�Myg����n|��1�[z�/��MG(�:`��u�[��:Z��5���.�ӎ%��w���i�G�y/ ���Ma�%ws�t�oa��ڀ#$��,o�D&/Y'd�����4��30��b�D?�w�_��k�&�Hh��?�(2�lր���s�.�	G�/S�H�跄�E	5En{�ҍ#���.��k'�1a*`@��:G7Zj�EմZHW_���Zp��LG��~=M��t_b톴Y7k�]�!��r���p�j�Z���z�o`Z��� d^�v��}� �1�J��{�1S��u��?[��.C3�	�����%��d)8����¾c~�mP����띘,9Ц��K_���B�><��t��Qט3u����F�����{�>��!��l���S+�o����]�8��Z�~�i)�H�[�۵�\�ae,��$�E䠅���ix{L�ɷU��<�d�)Z��Qx��̡`����MW%sO.9绂e|��t�N�$J��Oyp�Q���l�b�
;�0�Ż�|����W�I��	z�9+Ú�+�W���y�z���\l��� N�9���S�~H��-��G\H��kGBN0'B[�%(Ao�V��R�[i�p0gH��r:�����P�#wI=_/�<�+خC����u"�7>4#�� ط�a�ȶ�gpD�"<�Z�
�>�>�SA\z6-Ih��D�wL� o]BD!~l ~���&�ϻ�e-��pW� ����_�pM�8q-0�*�Ư� s�4?�*Lq�^c��-:M��R���F,i���'�����k62 ��B��6ybI�Z�&�Dy�n�4���&��\kѱHl
��]�͝�eE�g��^���i�땜����������XY	.3R�T
_����9q�80yˆ��`7V��1�#�Bx,��DG7��i�{Ym!�􀖼v�/�v~!?W�ײġ;s"7��l(�I�FnW�x�{�����;����e���-t����+�G?i�>L&���ζU�وOXq|c	���G�+���i����M��4#�К]bzj���l�Ej��E���N���)��:!��E؃k�鬩W�u�����˷���{��;(� 2�j�����عnJE��D}�B�q�恚�Y��%�?�y�/Ū�� �{�7�YG=6-�����(D���Ś$z�>��I��7^�=w��4%��|�A!������C
����ƣS���~�iw(��@�{�Nw��_D?�p�^�@�f�u3��U2�ܘ�#�ɧz�,�o�=���A�d�`�3��⦮�
��v���k�=��^�� ��kи׏aEx�;EDSo�s�'��^Y�͓uʶy�S�3�*+�<��b�o��-n퓗ѽ.�8�{7���%�|���J7�S�\���G#{�h�B��)��픂�L:#���腖$Z�F�Y�<c�A�J�w8� ��Cm٘���B�-�)F���.�sa���׌�y�^U�7����Ԍۮ�(h�L��:T�]����Q<�m�1b��۾wHЬH��b�
�Ɨ?<t遘<���g���?t��|7��+�䏿io;�}�%�=�t�Ϥ��Z���9[\�%�� @^�?v]�B��*�<�4���a���i�}2t�ߩmc-+�������N��dH�g\�K���=�����W��`]�eo��%|��Ͷ��N.2g��t��s�n�	+7U�[�U�t����A0�Ժ���c��n�;Vj��$�Ө���U%�!��Dl?P�l�Xj�\��+�͘�;T!Wd�4ډ&	���,u�Ųx���1���J�"�a��фn��6�3��XlxV64EB    fa00    25b0;{M�x����XF����������㧔oB[� �&���u���}g.�5s���K���:�K�I}���./���sƼ��V��`O�f���OK/	�#���	�r9s���"$@w���T�#��9t'���-��1�=�bo�?!ߕ3[D|�bSd��:�)��fa�p]
Z�G�7b�Y��~�7:�;%t�'_�=hަ+�_Hi~�@A;�R�|T���fDy�I�3��/��5�-��P�QT hG`bd�m�4K��ߛ�
tQ���̯V�vP,��N������˖B�"�h���+�2�j0���_ʵ;�X�z��?|3�leC�>�Y��f�����;c����'	�:#З���ǽct�e�����55;2��7� �kݓr��(Wy#�l�o�(z�Σ�c2v~�,̗��K��	I�IA�/g���� xdd�v����"'B�ap�v�rW�/��Q!��dw]'��֢�3���[�� �s��}�J�+�?;�ͱTz�C慨�����n�r���J4��hǢP�Q�C�ɚ�/Z�j'9�|�,�5���f<�����4l(������9��x;�/s�뚧b� �CHH��8u�����Q��n)Jш���c��V}�:�Ҳa\C�h���D�k�vm��a����#a�������"{U�8�x$i�%�~+t�wPo�[�G~p�T��׃�ͦlQ�D@�UA�<n�{�!���s"4�oaVz��5F)���R4�cy"�$i?�C\d8Ձ�vj��T{�b�����/f��_�U�g�
%P6�:Gْ���h�[��)20���y0`�gßt_�!����qG�V�%��F^�9><s���K�"�ݿR�2����^n~<lFl�����^2����q1�%C$��[�H���,ՠ����ɨAXhl�Q��U��}8A$s�E����p�'�����)�g��
�(lc���8��{ת8f�vj��V�5D^Q���ÊZQ[%(!Pct��\�Ym@:�.$x�/���Hx�\E�l�5R������t:T�@)PDdZ���"���zN3n�U=j`x��iT�UK���"�(���I�p��cP�HGکA[~����޼'��R8�0 ���h}�����+����r�%�N��r]!ZCK�~Ϳ�����^�:���c�I����R��ksk�oo�����/u���*��+ˍ���N�Wu��-6o�����CT��MӝѰJ��#o�u��u&C����K�,Z�zS)���Z$��?ۀQ29q��>����jWS�0���ˡ���d�U�9PϬ�>}
�?�k\.���Y�\��5�������q���׻ϗܤ�2��C�Fo��Z��Xl��C��$TB�8�����{�Q
��\6R���Z/g�"Y3U`.j^E�4�<���`��>�cÌ �����Ԕ+�!Y�r��v(uK̀|v[[״֤?,�Z>�,�}�$����}3W����VyYQJ.�Śv=[L�6�a���F���{O��;���2�x�Zd�!�wd\��~>H�?/�UH`w�< ��*L{�A��� 0��5�b3�`���eB�K�`���y;�o[h�A����
,0��5�u|���2������DQ��FR��9��3o��Nz�`�w�3�F�n�9�kVA,��f�P���Y���S��Έ��a	+ۻ��n��Z4&���8q}+�����o`#^p��z�>6�[��%;�dج���X8�E*d�5V�,��� ��5ui5#���iޟ��!u�l�����2�y�>*�~^�r]BK�{*Ӛ�ra����(���g~�O{�b�|������(Ekw�G۵ȈB��p�FB��D��}V>;��EΏ�7h�|7L���.��܆UNN��䇛T1 X|~���S�ߚ�� �=���4�n���,_�
�.Gi]��ՎiUQL�8�#&ӧ�ĸ�G�~�D�(1���-���x�vҔn�T����uE����9��n���X&(���xޗ��s����l�e����.�������y��OR,c׊B9�e����0�~i���3��h�\Z	5��布�K���������d6`9ݿ�{Ӗ!nϕH3��s�
/*��3����X��}Ӑ�Dٿ�풣4�MP?��-�^E�����1���՞�z�-'��<���?�]v���dF�K��p��;ES��?�S�:Zh�ϭ�V]��7� I��u\�2�b� �3�_ ����4sK���h�G϶4��ɠj�q�+�G	���� #?@q��jz��E�d](��m���S�B]k����{���2<N�y{�d� CQ#���k.�w]AH��SVof�9��]
%TK!c����6����Daj�`���s]��MuT"��q�h��Ɖ�`��'��$�.�|�޻�.�/�����+�-O� 9�J�U��Z�l>��f�h��U����Y����]�ob��ZN�K�H�/��l	��7� �h�Xu$I�B�Yc:��ɵi�}aMS�J�NW��X��uo�*��1�"H��UlS+�J2�82�2�j���Hu{���p�Y�
���P�0mCQ��_���-�I�t�Q~��oC�t��"��\�!x�4z�a�y3%�I&�uVq���T��n�?�P��X�̎�
��h��B���z�_���s�Ay��0�������|��?�j�(O�!���ݷ3�Z�Hڍ/ד��bg~��IP	/�?��+L�ތ�TZν�[�%�lPMceݑ�q��8��!"��-�E@]�<���]�=�;�g�*�l��=���f�wS��n$��q��8z�����iϘ�\�Ow3̆xvkr+�~ξ��ۅ�J�����e7vݹ�s�:�a�����)�e)�0>4l�z2蹃��w����b�r�Vh�Z\@�>��@�z��W\��3m�a�F)'�F���L2��,�nf���]+��G�1����3Tb��G�8��x��2x>������Hb������)�z��%=��bD63�Nk�ثT�P�`��	c���z~V���F<7�$t��R�M��M[�5����@�N�pP*�N�����aŶΡmtf�ȹ9o�n�F<Sp��]����8��)��OI1� ��Q{H7�[f��b��Ϣ	8����oq'2O�w{ʩ�itk1�r24Hİ��m`k??�T�i��ƠqT���I�Ky�����x
PI)��8g	Gz�d��d��K�m�c������L���h�|A>9�P��2�l��\C,��C���9�dRemzd\Zj!~Xť�H�;ҫ�Z�r&a�!��/D�1�|�C8�og�:��t����ԪR�%]:��\p�.�9H?�r���7e7|F��&?&�� �,��^D�j,��`�j �� ��Uu�v
']4�LBUU���T�{Dv�3��`gH�
��U�9�O&7�4�#`;S0��M�M(�![^��[�p�ձK�s`f�����j{>i�ƅ������^�k��k�Us�!�:T���<�/B[
vF?!B3L���?[�� ?A�v7fxm
��O�Ds�85��xE����z]`�+�Z�, !�LC��3�����UJLX�՟�-Ʉ1���j�GC���ɫA�����^������M*��o��*��F��ɕw���%j~@c�����\�=�g���3_�F���cȘ�0�oVy�4(U��2�!�!4��2y�������wzW�j��H�LM2�W-�C;Mv���5�:
�J��7R'4zÒ-������	��Y�pn3��[����7DB�.�.}^F�%�<5�S�~�.V�A�)7��\p��/�r�7ig!��!��;�=����آ������V�`�`�I�j5�a�IL,���$�tc�B���m(r�5W�?�����s�l����u2Ӵ���v8����m�^Q��.�=���s����܋��W�����ԕK���S#J�w#F��4����)&D���s���zu��s�
�l�׀YU�:v��H`^{�fQ j�5,�
�@����5��X[M��w�BK�Z�U��y�Sһ{�/��c6r����Ъk��v$UY�P�`��YlE(�"3��5;��3"�=�]�4b�k,e��[�F,A�e���^{,ѺDpQ�����L~��1��$�������^��ی���զTI&�|#�B�5"�f��'y���^d9V�x��聳�-J�+
\�.v� {�Ċ���5X�l ���B��iz���q�c�.eV:{�XDh�2L�Y5��F0B��#�Ҁ�P��~��{d�Hc;����ζ�O�W�Ǌ�Z� ���[�W�����9��E�#��A��X�#X��_�,�`U6�9y��e8���yi+��X�E�o�QP�f�T��wi�B����$` ����-N
X �>���|��?��؃�\����U=O��TQ������h� �W"r~8é��#��mmh����n���94!���A�W�A욝/�Rɏedӓ�FF��? m� "�q����UI4�O�z���k�l5���y���0�2�����yH��i(�w��Y�3�]�\�2�@.�?/&��q3�p ��]����s�ڳ<��'��>J�l X�mps'�{c|��������v����&Q�����T��������M�Y�U�M|��%�1�A��ֺ�ڍҲ�SE���@*��Ru*�e�z���D�B��=|��7�l5sN�oj��R4>��&xI��$�	�"~����!6��U8�>E���|Q�������Zg��l3:I8eT���}W�a=��l��k)|+�%
�♈���l����+5\�a]�j��Q�(#�Q�c_��b�㦉�Ʉ����=y+�!��[G{|@�g,�L �ܓ�����Ah�#�&�@T3�.V��j��h�HS��A����%�R؀Ng�՟��!ㇲ�}JͶ�����Hd�*�4��zBvaX#�|���S3<��n�w���c��s(�~�>!��c�}��4B�殃j��J��2�z��SB�i(�Q����P'�xF���C�U=c������۫�fÑ쐎E(��DXmhq��(Z/��r�N��3xƿ��I0ߌ�$��{$��[3z�Q�c���P��4*PO%�D�S�7F`�:���I1�nm_FTY�ɜ�u=��b\G�t�U��O�Ur��z���XA��<R��P�Œ�ɩD"���!Q�����/�u�}i}1l�x�d�)�j�+��f��c���ܧ���#rn���_h��e$E�l���i91�O���5���e|]�P
)��e
�צI
1�#0�DZ�y�s	�a���U�K}"�~��|�%�X(���Y�R��S�5o���lN��L�#�ߡt��u�i��2�t��$4�'���^�����Cjг:�H;sF���[�A
|v�m�3!b=x���կ���ܑȸ)nXi�.�� {m������~ǟ�y�g�w���)�u4�W���1~��͑s� ʷ�@4��j��K/�ԺP�y���7��o4�,:3��23�j�,���L0�;_#B�N�!�w�-��c+���,eR�7��&�O������.I������X�WQ���~���mu�/���'�����([��^�����oByjv{�C�A����:�_��F$���@�!�1�Z��͵����b@�2���Џ�L�9`�ǉ�بжH�f[�z@�{�"gY����>���ɔ���8�[��G(�����%�~i K�f�7p�R�Hh7��O �s$)����t���0�ŢlWnO5ry�%pF���>߂QJ���9o��_��#�VA�D���\:Ԏ��E�����+�U1ߙ�j ��N�5;��Θ���@�%�q9�ih~��d[�tt��6o�[���1���L����)��?K&�o�
}����"9��_kb�s�!��S	�����߻��~��>�#'9��x��xZY�i�A����@W��=�_���wȻ1�`�3��0��p���D�H�+
+�&Bnw�l�,0qB;'�`r�P98�G���n�,$NZ&}�O�O_ߜ�$� [o�����P�,F��l+'V�����K�e�U�R��cijVw�,0�rP�
GN��I���g��V��J��E���M=��b�����"�N�*�Z��s�t��^h�	W��H�)�ێ�����o�ɺE)P	���|����N^�01�.��?��Y���M�|��ri �g�`���icJPd/c`\��P����qV��ŀN�٫��@�3$H�0�=D�]�	E�l��M���(��������E��[�{�7��N�&(�/`59�E62de�6��*߸��T�ʉo�÷�l]>(P�b�$_EU�E�-	$�:������\^5�)65��z��KYS\�]րфn3��X捭(e��T��J�0+ʞUz��=�.�;�_z�T��0V(��xLoX��h+��hg~��N��kk��&3� �A1y�~��	*�V<T����{k�.���[7�{^��R��u��1;���,B�3o7�X��4b�6(:�򔷛ݛ9�u��!"��տ��
�j�g!Tڵp�\ayT����	>N8���Q�g���3A�#P�ͮQA�.E��C
�ʮ�8��a�_\Y���d��4gA�|��]��D���R��ìD�дr���5��IN���ɾ��R��o�s�F��k�č$�(J�h�oQ�!��J�<q���\�+��� ]�Ҝ2	����@
����_T������-va�������R�Y��/�l��Z�Ӻ���P�̐J�U�l�a���nI�Z���J��i�A��`� �:'������d�J*�8��<p�5<W��8���~�.�	>� ��
�c�]I)�3^[f�;�=#�q=@�%y$-���7�b54��p��c�E��Z����=7���A2o)�t*x����,�"�w�����th�ݤ>�',!
3Lfg�����:,�S��g13�$�S�q��u%�����ئȐ�B��Z<f��1ߠﯴ���В��U56b�]�9y���9T�Ş3�;�^8�ys�D	rk��I�v����@Kj&�[G�؏%�b`s�x�Z��Q���dPl٥��"4w�)3%g͍g�(�im+��5k�� �3[��'fa�Ic�� T?k��p"��wbN�%)���nh�sİ���y�3�j�{{�W���Z�j=�M�bg�'�qt��b�3���=�TS���o8�b������9�F�3`����k��*�3N��a�R��e�Ͽ�C�%��UCz��=/��l���G���$Z��z��ə	���Z3���ڲ!���ɢ`W%����¼_y�_ ����=q,�6Э=]�5���N��q�AxXC�U�5U���L����n޲g:0�j�Et�@�ä�V�Fl`I���tC듕�A�h*�q��NhN%i!��ͧ(d�u��X93ή�T�!����8Z���
�/ȟx[�<J�J$2G���4]4�� .OΔ_�:���!LF��s���~q�8WH���Q潒�''�Q�ˊB�ݩ�ޜ�C�p�F���[�`?5|Rb����qd�<H�2��,��;,�o϶W���L"���LҦ�y!�B�a!���kjb�1������߳mL�uG���T��"3�*'��Y��)D�x��E�P���qN_YT7-֓�a �@���#��HX\V,f�B��p���l�Si��y�':�UdB�Z����o�oL�*?���屷�X���p膠���p()��_�Ⱥ�L�\�T����c��Sc���nV�(������X��W������>P��%{K� ��獳A�֝P,�M
�N)qJ=�L3h�z�$?ě� �\�P�e���ѡ�(�75r��1�#��7{;رi�z��gr�c/*6��ؕ��VH�����@�rS8�C��\*|��w_XBj��s�h>Hf�u���0	|	[A�~]��9��N�I�A�w�w��}r�u��X2c�qu����!:�؃
�槌C���O�	,�`#Ȧ����.$���<{}P�]%}S���}n��i���I�*���:�AA�1��H��t��(T����`y��X�L�2�k�� �(9B���2FB���R���G���M�|�_�7��UF��ϑ� ���P׸0d�.l�6�=C닶�F��<}D��w��B]@���:�'�#b�H�n��,N.��q�����$>�Y�\��s�"k����A�vo���vTli-B�,Ͱ�Vջ��ލ$ZO	�.vt��'��IV����j/�	xn��d��s<��m�`y�И� ���/8�%�"�¨$S1޳N����r�s�_���N���	w�[�Z�!z��_���5=��5b��͝��+ߙ��0�=*��?w���n+h�=�{��w8Y�{�Ua�V�-�=*�4���۬����*�����gh�r�olY�u��7�%�vׄ荰o<XR�u���������Ը!��6EC=!�:��/(�$Z��6a�]ڌme��21��
Xy`�[�ȋ��E3�kj�x��WJ֐�_8z��S��`����G�:1*)|�f�A��m�<�
�s��l�Сg[����MG���|w��z8怆e������m �;���,1+2�4v���{����0x_F
vg�K�e��[���	��FYKt2⛣����m-OO8?�L��*���a� Yu��4��﹖����W�S��C�∃�\\�q��@u�e5��q;$Ŕ�E9GkLV����/7󀨄T���Y���x��.�����.=�B�,0;��=J[�R�JW`�UT��it/��NE�ho�%~Si<A�t�H[$�� !��ȍBmLy�TW���';z�(��+*S�x��{�!�F��������Ne��i>�z�N.�(0����'�"�?�{�=�D�	dN c%$	�D�5��֮3Bn7��7]i�Nd���!X !�~V��-`.��������wΦr�]/�@�S���*�X3`Z\s����NZ.���	-�W�������{��Ԯz��4�M?��V�M�%����X,�\�ȷ�?��0���mb�2h�gV�����Y�{���}�Ec$��1���`��I^I��V+��`����<���\+5�F[w�' x�����Gu�S�ꛯ��b�g>s/�]��q��D-�����T���.R��\��¼J$\1�\ܛ���������"��߾�s:Ԧ)#!aF��>31��I���q�%��s^C�ݙE��^�q=gyZ���F�,��?����-�BYt>�V�s~~'<��v�g��DM�
Q���<&�k=���*��bZ��{E|�Q�{U�:s2������jP���y��K[�_6��R��"}���q�ױ�~�!pE�j/��XlxV64EB    99b3    19e0�!� ��vMu�����_�tV&�.���j)$�r�x*ИK*6j��G�����i(�W%oh)�}����V�E�l�S���|az�
�{�}�c��g�gj�!�Ċ8�V�R�S��)F�i?d��_��&�5�=���Ǽ`�d#dR�a�I�K�H@�G�>�NLƼ�%5�4�Ο�\�w���ұ���o�s�Ӵc�E1d�p7h|4��H�����O\�b0V^��s,#Y��$���KVVL��8�&�c�@����M�ǖ���h>�R�73�2@���� %x)I��?4k�f�;��t�|���Y:����s�dp���`��TZ�4����J$[:�Y%���A-���-��X-�%��������B�:�ݯ&��jwM4!8yM��O*W&!�wVw�N�BV᝚d�B�?Js,�mv*�FmC���L�{a�R��	Ls=�'wj�oP+ɢ(�[( �~�[�102��OAj�@�Qw��$�t?�n�m�ql;�17�'0�]���l��]�8$���ů\�A:�_ϭ�d[	�iK��e<������'p&/�z��:ג�=�^�� ����\�ƙ`v�6��w~Kd���d��IcL�SNX.��cð�.�"�BSrŁ`Tqr9pf���8	��<�	����G�nA���|�H�J-���֖�R���_�>Ͻ�S�MAEvP��>Rʎ�R���;&
<��%�/�0o�`1�P�]���D�.  �G�/����-_F{BË�"��(�kූ������I(iXswX��p���y9��u}~��}�o��s��|(W�����1�+痠���D�p�3�(��uu��W'χr������|Y�$'1(�/5M�$�Gr��-V���#�2w݁����H��wx�CɊ��٥Tr����/�Ur��d�5�Ն�Xu��B���^H�l"&Bӻ�������H6��4dX�V�VF�}Mk��_B��A�}�)M/ǡ�@�aD+���_{m�V�0���J@� Τ&��[��p:����O�S���!��_�����|~@W&~��v���ҿ��/�'~�^1�ȏu�:�!�(�}�i���{��"���D����u���ks�2x�L�.G�i�l~K+ބ��~��11�ʆ�|�4r���u�Q�1�V.��a���D��9�����G���\ X#���ۛ�N��@P���"J^�~�r ܞs�wz=�[=���_��So��+Us���.�ܬj��MKy%����C�B�K�����}���[U5ugu=��j��F��2����^�;(4�[L/�ɃbӐ�+�KP����P!E^��̒��2�<��c���`�PJD�&�y�s�z�WW ��R�%���ڂ#VuG��;����x����Ɠ�b#@�!p)=��*�L�x,4�3Sp���cn�r��	��wE��a�^MEԻ(*����7��ɾsyӹb����o��Ć'f0nց��/���E((*�Z�m$C��7�m�A�d�l�Gѝt����m��7�����Fm�S��e4�N��m��a���)Cݮ�0�4�	v������op�=>��?�)'Sѡk���Kd�G��˯���γo=y��Z�I�������<"�놠�e)sq�-���#�(D6������@�H0&������J��A0������ {L�F�e��Ir,�k�Ϲr���G�����`��d���6����j�j�����(���o0A���5;��|+�?Mc����`��,�mkF直_y�-B9�oT���vvK����&�ùh���r���HZKn���g�Ǝ�+���Nl�4+��U<�J$dC��a��*S_�k� �Ƈ9��q����	v�%�LI~�^SєO�
7��e	�g?����-�?6ڝ��v���H̋����,9:B �4NQH>3��(��!¥��4���Z~�~�)e��g��}���ƈm�	'�W���n>]V9&l~Ɣ���2n�?Dg��i�T^E�#]�I`)8>��Tg�_�٭����Mu�L��
y%*�E�L�4�ѡ�����5���N!�^ą2�~a1mv�sT����b�x��k�'6�O����P(3%������,�{�bb-��JB��7iFav�G�f~b�[TA�s"��/��|� ���?M��Wk���v�����^�Z��@���nJ��ͫ�yYD�E}����G�����_����%��/"*a�J�K��PClMrwm;H��<!4_�W�}.��K oq>�M�����f�����{�yWƌ�{ɮ� .\��Ê�ez3s��>� ���8Ur��W&�0� 񙩺e��`{H6���Q�r䢋��{cq��yv�qc�p������K;��F�G��r)D�uI����������iK�MW�"6�|䪐�΀�4 ]4*zv�D3�o��Q���'v@u�I�էC��qpg{��V��$O�Ė�k<�$#�)��u�"Y���./=��>S΄ �#Er�-X�c^8�S�X��#%�k��*�x������@�#a؀K�Q� B�L�W,ͨDuKsI��u�e��k�4��rv=�C�lo���Bj�T+U�V 5+ �Fy���d������ԋ���id[n��'��j���4�W����ЭT�N,5����tV������� ��2��lg@@A�� ��5f2�s9�����f�v ެ9��g
�ߍJÑIɲb���b�0��$^��档��@�q���k�����YR[�nn&��"�'/=2��٫��0����P�9�i���N��촐���i��]5e�t��6T�Z0ZE��^�?��(���}k
N� X��nC����1�O詉Y��Q�M��`�TZ7ڈ�s�{�J|�����[�?�2��Dj��kGgI��;�ؓX(��e"�7f�����>09��������i���볾�gM����r�}�
J)5��TT�V��j ƘoM�w x�����n��(�ڣ��l����ż�)�Ƿq8�N���Ê�V=e̅��]ݠ��潾�+ލ����#�D��1�����>�a�9�&wq�
�Ǔ��syW�F��:�)B���mU)k�oji��u=rqPT��FFhee����Aq0o���GS�����qkؚ�����O����/0n��1E��Ӵ��	ZL�_��,Ŭ{(,��H��+���Qڨ:��|�X����J	� ���2�L��v�LL�*̀d�~�`��F�_JE�|0�V���3�F��t��#��Rey���Vcew=m�<���a|hì�gu��u� ���x�M��B�2�`"�ӷ�L�p`�yqV��&X7��D6�
���n�_.��ϑ�E�.>���uy��ssG����11ݻۆ,�RhK����Y)�5�(��U�����ͻ�'�q H��J�2",'����?�� �0:����;8P���N�^�j2����nW̞��BYh&�ِ��$�0�;�~3��b�
G�� ������蓘�p�ߢ��(�xt�����GS���l�&���g$Dx^ވ��5`�H�i'``	ؼ\���(���_�ϻ��t��^6� A���AB���g�z ���,5b}��s�
�����m�k4��رr�ۋ��G�5"rz��X��{�#�f{�ʶ�Z6�:�3����Թا��1�np��!y"���o�L���_\�AL��r?K�J&�`�Z�c�`��Į?�}��+'#�3�Fd8��y\��&r�Z�&^�60�r@fӑ6b��Lg���_Vc(�^J��w�-���^<,Ê�r5&^���;�@Y�I�OR��w��U��O���H��0I�a�3B��*�'L=��=��@"�jE})U�x���@��B��U��
����ս��C�J�"-��AR!w�ea���=υ�N��)�O���;2�]�z�7V��_L�+
�k���z�"��~��\i�>2 \�C<�E��s	E0��ƾ���c�(�F����q�Ǆ�`�BJ���xVB7@&�I�;��+���Ѷ���w�9�@��y۪���������^V3��z'ը;�k� 0�o3^�Zwp/;S����߀�b˛K�+�n2�Ļ���楏O_xX�۔*[q�1��7܌�)t�ق4%I<]����kK]�9�>I�>�"m�P����7��RO�J��O�@����?�ܟ���7����Q:�.Eu"�!Ê�2�n���j�'$������%���4ұ�Z�T�2"+#��qJu��t�|��!N����qM�/�5�����z���������(��,}-	�̎6�XP4t�#p�d��[���[�N�<��^��,��u���Z�S�,gQzꭗT�������V.1��'�Є&0�c�{ڈ� u�U�h�A��#x�]L��Nn��g7��������$S��,�OJ\ �sv�DJ��G�����d:���g�s�=�rl�\����@ƙz l��;�Vǰ^�:�:U��Q�`|R�*mH4�1����r.D-k�n 5��h�CE�y�	�Ф�i��e`���!�ݼ)�d����r_7��]���($�g~ș�t+p��w-o�#1�3�.C�M[c�7�8��� ,��X���nW	��k�P�7���*�lEَJ�%H�	~7�2�i��̍�է+����O�����2�BQ�NQ�P! �~Q�S��HK֩'��h�G��ϖ�'��ڭ�=='j��F��s��Wj��88�n�{�9K�����\��Wz� �JG�*�;�z���J��v�}���G���������ɖ;b�a��ܗ�P���u���ϾŹ0bЎ19�����'�6�kir �'��w�W��:�yQ���\�Db��	:��SP�L����'�`%��(h_��R/P�a�{Z�������E�6�|���!#����g��ƶ�&{��p�Mh��R�~G��֚X8�)�Z<ֻ���`9���P�� '�U䋞ڟ�-�ߵ�t�>\,4�bT�zxJ[����� (���)c�t���� 5�V��Z���R: ��|�Muj�C���#j�e�(�w�3ǼƄ���/�`U�/-��C�=���u5�4��]�,L�mɲ�hM�cP����c�Ӣ����������O zP���$W���q���� 1#�z1��7֨�pV�+�;����=/;��)_t�#��'�W	���g9ǌ�q��Ȍ�F�b08͐V�1�9��P�zf����C;{���UX�zkDy���s�$������ w�ҍu'[ҧb��ޚ%K(<=?���j��Z^n�s��*�Pp�0��F�S�y�o���j.�K1B�9Ͱ������غ�e��b�?�0�g0��l��tb��;�C�DLj#�hȥ���!��.3��H�g$PmOh#�V�{]n��hp�$7�IV$����q�p�'�#ag����QM5³m�K�٧;�Q^O�H�B�K�Ъ�~z&�L�뢻�^��W=�i�n�VOM�s����D'���o�A��.��Ѽ鷻wB)A����w_n�em9�"�B����Z/Æ\�nD/q�)���c��A�\3P������,!3"�*Iׂ�\X��&�wv{FѣFį��!��-3�?M�]F���q\�q].�0�	z�O�%I[RVo�<]Ɩ[l욱(�����H�Pƽ[Ώ��m%���E?��p<�8��}9��}�D�`�� Y�#��Ċ�F[�F �]٦��:�I���9
p��&��O'%�Z��gf���b��?O��;�NF�0b.�\����lIu�$w��&�=��b��$�*W�	g���[���fj�3�Y���dH�-�\��V�0<@�T�M��oh<QbZ6��q讧���D/��FhY?8[/x���U�Xu�f["�=��PJr�`3�=���t��ۼ�Е�ƿD��3/L�*a��A�"�_�C�Y�����7D���4K��yzP1����|�_���(�8���R�R�n���EZֈ�AԻ$č���fZ�!�(�V���o�=k�����:M�j�t]�#�5b`{ �:�Ms�ZO�����{>4pc�����)�5�O�Z��v4Qa}����$����KΌm�v� ��L��+tY8������H���Ufuf�S���:sx�E���sm��B��S&G��jV�_Z�p���7@�6C�+J%=��OƘ�cՒ�t��ܾbY�ʷ��\�� �G���g��ϗ�*7 Ji0��mJ2���A
�M}c@Z����K�D�oh���*�Z-�ⵛ��y=��� 4�ue�\�>8m��H�O�s6eU �V{hjy��6a�E��u���������b@����^k��L����Ah��s$�5��ZƈKKx�~U�䈞�e��!��R��KzȻPcS��%�,�O6I=�n��Ҋ�Uw٣�P��y�= QN�J