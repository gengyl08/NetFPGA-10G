XlxV64EB    fa00    2e80�l�W�I}a56��QG]
�w%��z��)k�0�����Ƹ])�s�\�}F	����Y�I�b�̹�dխƆw���̆;��w�L���_�*�
z`��=ۅ̵�`~]I2�z�������d�C�!�'�Iz$ �q�i&a���vb���g9?�u�i��%6' Vm�ٌ�
bpz�g����*�z�&��I��+�r�]k,�@<�u.�ѵ�鯽��� 3X���=	�ޯb��t.���E�h;B?�j!�O�&-O���$R������z��l c#�d0����$v2���,E�È�\f:���)m��Bԭ�7N�
�ܖ.�̚�f�=�fk<�̎ |v:�BybV$a�[�'�z*�������ZuE��a�4��){d6k@p��`W�����~�G?�]m�3��!�HL;��(���b=b��oY�?�$hA�bG�)6�w�`
��}SM�����ٌ�ND�6�4�v"�PY��:���5,5_������W�7�_�)`��&��Rq4�)KI��8�Dv�ꚜ�r���ρ���EU�S,���T;�&z�ǵf�h����x��C�k�@�qWQ�����m��� �/�e,��=�|� ��S�t<�?�cF��D²EڿNF�W���RN�o1����{�^E��Z��� �2����ROOy܆tQ����V�ZxJ�?]>4.f��6Am�L�+Hz��?�m�M��#���x�"�~��2�	)�}$�hpÕ��zc��+��ji3C������E�~U��)W�9=v$V��q5n(�6��+L�:�[آŧ-��>�x*L�Z�M�	��g��S���+D��ZrI#{-;��`�h#x<3Kbo��2F��=�Y���8#���Pm����+CͬfQ���z�;�gx�7~��h���+t��[ք�V%Q2�5�q��E��;Ya�(8x�ڈ����_S�ɱ�<oHOQI+0 ��e�����w�t�c�;����C�֪	��' ��Ӕ�3��n�9I���q�1�A��S�@�|�$&�K�ȁ�n���ne��D��%�����E�q���拄ox��v[�2��b�ĥ��*C��)��q /�Q���'|B�Q�R�M�<���=�8��~.*TDGGb2���������!5�@�l����\S,�����7:&Lmϳ�t��ܛ�E�s����3�l[x<�_�XT���_��o�'ߕ��QZ�_^8j��i���3Vt��}���h�;�W�>D����B����U��+��H��P��MQ��jq�kw����/�����uڈ@�a��1�4xXg�����n��U~�3.���i�V�8o-խY��K�G���5�[���S��-��}��e�!Gg��k�����C=�������ҁ��p�?���%6���#���R�?�s�k%JN?��)NNOD4�'F��o���A��٭��<#��7���y���V�L= ���$=�*�qMKFA��5�ΐ~��8��D�5��P�G�<^�F�r㨒?S�R�cK�u���S'���$[߰u�@����M[Jo4#��2[	V��m��m��
u�xG��t0Ύ�e@�]~q��|� N�>%"�Y�%+O�:��V�?ߵ1�,��ez�/�*I�����{��ű��P,�] 1�����٪W/�����d��պ��rqd��0�l%|V{Z��?Z���8���O�x��b5ެ��d����!M���/;�}{;�&�d��k�A�:�Ehv�V�ឌ��SU���sªL�Y�h΀�]8wԡ�6,+�vכ�����Zl]t,r����ND��2�8?�h}f��O>Ů:�
�i>�re��AY�}��OG�Tɭ̴Yy�8��� ƹ]�c+��'A���l����U�1���@-~�)]_��,Ч� K�Z�x���)W�I��0�
U��q�]����|�0h�VǠ%��^�z�3��g^���(r�w��֚1O�G����^u��֪���-�ՑX��!�ɮ�Z0�H@�M7e�����F�_��7�ba~֬���p枃@5�/˰��ACIۤ�ZK��V(����[�'�$�Xk�Aյ^k�z���rp�K��n:��/�Z��-;s!�Z�Q�w^�������d�R�V�V$na�<`�xފ�e�� �n��3B�K��Ҥ?;q�x���<+���i�9y_��� Ȳf�b;��F篲��'V^�MM�/m���RXW�r��:)��(l��`�)Ľ̆��-qY��zML�ޮUNu��%�"ٖ/���*Cⴑ�m�ģ�x������]�FT�O�?���Y�[;Y�7�ݘ;� �S�m�b^��]k \��e�r�V�gry��b�F�nb9��I��qm. ���6{C�[8[�9�%�_�Q�e����8�#Kh&��#h�v"�@��I{m������٪Q32��w�j�S�ǄԭK;� y">����J񰚴Ǹj�x�.�B�.��`(�;�cf
'c�phJq�3+sc �ޛ�EWE�HB��u��V *y�OC���`y�c[��ɇG��#O�;^�%tC��,�QpS��/���w��|��-�����w���Uuڛh{��	ڥX�����c�¯�,:ÿ]��B�=D���]�s����_]��ѱ�&�,F���׍�;�I�U"IՔ�EiO�O�Y( ��*��G5��a��6��'�����Ԗʗd{L���$cvX�I���"��.��^�CGl�p�l�WѠ��o����\��I~h'S)&�M&��@ھ��H�B�5�g�Y�qǬ��OeיU���ho�A(�˖w�Mg4;aʵ�fY>������a����m�!�:i<���g�Al�7���-�����I��{b�q��^k�G��	A���U�h�g�iW����W"FQ�Z�ŕz�������K0p�4o��$ae�T6`|�k�0*:Q�٦���6�`p,0���G*�4 ���>[�a�(��G1!h"��=�#�-\}����/���y�~�_?"�ȴTO��{�\�����q��0d &���¨N��Ri�5���o]!)��'��ү��F�����Xr��5-7N�'jp�:<��)�/<��^
�Mhf���pF%�2�z��p�� �)��������l�%���_T?>��`Vq�:�%�2S��)�{����14(�1�������I��f ��a�_#��ڍ��m������X�ؿ�Ʌ�� tr��ԏ���s.vF{HN��6�e���xi���N����,����4�R!�[
A���G������!"�u�x�LnV���TaD]Y�?A�,���B�{O%eG���n��B�u��STA��-(�P0�zɱ���*������G9S��b�y�.諠�y�(�Yf�f�>�N
:�hu%�Ul2����Dܧ��Z����%�dF�#1������d��xe��l�U�b��K5���K�<��w'3SQœ�мݔsz�V3��d���2��(�!jv�W�&���T|��DH�����9�n^}��f�۴/ۤ�B:$D����d��ߡv�L��B��Ũ[:��F5쯠�$�ܕ�/�]N����+Z���2�S�k`���6ryE[	e�����[}B�0�\��Hj�ۺ=��w�)��D�k~�K����@^�%<����YBݜ�6+ͥ��%��/���[L>A���CD���� ���y�zw��]�r�]���f�w+�� 
 FuO�.3]p�g�2��W���"^|F;���R�j�DЌ�;�8��/D,X��O���Lk.n�C{����{��¼�RC��wRgji�D]��Y�/N8���������t�T��"`�4��d� o�W���(�@+G�\�L;�5C�}�'1s&����ygN�cn'�]�J$:�� ���x�z'����A���r����I%��q�fC�5����ֈ���	���{�ȿr;I_���;"57�\ݏ��������x�u�@%�Ә��ӆ�h:�Y�����S�E!�&§�>�2a�"��eZ�GZ�ӭqj-��Ԯ�S}�or^R֜ |T��q�D�g4$T2L�l��꘤���<��%M^qgOY���cm�ϕ���>��v�,<xȭ��䩇.S��'��ê�k�����4g�p�Y]$�D�{���=�<�?U>�����&���q�O��c$O��������1X�-�^��*�8�w?U�ќ8�D�"
�1dD��8p���ř2Y��6��^
��RC��m�P��8�i3���K���5X����Z���_ 4�G�N��O�ؗ�;�SB�\����J�γ'�,'ۀ�B��t9���m�tq/����?Ls)�gg�<���!,�N:R����v��j��j�������ˇe�x?ri��<R���w��@�Wc'cD��� ����}�`%�'�;F�O&�N��,��@�e�2�J_�k0�& kO?�g;�MB�1+��I�V0C� �H~L�׎�\G�@�C|=�~Th�E�7/-`��4.W :=��w���+��z=������K��>0��S�4���l���L�=���I�t�fWM%G4�m��unP�XM�Uv�2;� N���Q�����J,R�e���l'F7dh��޽�A�� ����;tUt�2i��Щ�C^���fJ!�[�~��"�f�����B�I@�;M��.6R�և�_�(4i'^�p�G�������Gz:���q��9�U����X`]�n �p�t�|3�u�i��x�"C��F�F1�9<U�uJV�Pθ��\�ECC��D�r���eq��U#�`}�h.�dE�j_��@N�����n��܏s=�Y�#���{�,V����Lj��@w�Ny���i �?���drU�/tz=	��rYg�k*�6b���'�.`7��*!��̚#�������!��Sl��@w^
��O#���D��M6�R9 �8�Vmf��Z���ɸ�j�FފZ��hX�b��n(�5+���3��4�8��UqE�p��o�c�LxVЖ�W���&t�X�g�0{v/���ʄik�7��af�HR$�ք3M�SH��M"H^�+ )��dE*\�VMع���N¤p���yXfR�A��hOG�*��A��ۖI/䉥;B)�l����CZ!%Rki�0�eaj'���OK0��S�j�#YnC6��[Mf�H�X�l�I��}��8�·t���˸bm'��[��k��`.��X�c1��V�SV@�,F/��B��v#\T61�Wq-)����A�8�wh��$s�%�	&,6�ҫxF�#�c�}��-�O��҈<?��3�U��|%�+�yY��k`�0��ӷҏ�D�%Y=���ZM�@��'��*A�6?�/7hÛßAq�[38�"u]֛_��;�n� �/H�j� Ж��X"��?-/jr�1u����
����9�����5{j���o��E�0�@��n5�A��k�Z]wEl
&����$|�����&PO��
�CIԔ�/l��d㻷�z�|T�k�j���`i����n'e��f38v|d�jy�ȶ�N�pl��kIU>�jm���Y6��� q~cw�"H��<�����S2�^wb����As��H�T�`�A�|��=�X��@�Π$k�����>o�Ԝ���H�P�'���A'��l̠�R�@�d}Sи{�����lr�q�a�E��w���R%���\��"�6�<7NX#EW�iE��4J���Σ��$A��q�q���9L�}�L�ö�������S�'
lXFQ�:�9(o��x������;�DL}f���X����y�o�= ��ڒ�%_��^��;��n._�H�&�M�{���n��|�����u�y����yx�/��0����oo9J��t�r8�����'*�Ŧdqr0��P�bݳ���K��h�>Rˈ�	��9TBʶ�����S�
O~���H�Z���g�J���3�ߖ�-(�`S��$�Ҟ�g����!r��q:[�&ǶiSf�7����\?�y��Л�7��G�3d��C�
�+ ��%T烥��b]���G�����Y���wc�)�\U�4
 �� �q��Vh̍�ܟp(t��
~��ݵ����/?�ײ���}��<}8�\ߣa���~Մp�p�zlP;���#f��9�X��5Qg"�p�G��-��q{�m^?����Is��p���'w��V�@�[Ӕ����u���8ߩ<$ĕ�8� NKu��41
��2�1>G�%]�Z�)[������O�.�Y�h����h�u��׀,`8p�hq��\�o���������(���j�vm/7��^�`�N#��Z���X<����1��1W�� cx��ًIzQ|��!�������샗����6�pW��Q��u�z�����?/n�������4����Z��S������SۊndEW��m���~p �U>�B?w97��r�؟,���5�f�eԦVʼ�J��ΐ�}��**�Cb����0�27� G�5^T�@_m��ɱX�GE��#���Y���#�Dzm>X�ڟ�iu/eR���BN��EXm�?�,��&1CbJ`�i��`����ų�kf���Q�Ӈx-1�;����J�A�B^ ��x���l����G3#q�Ȅ#�F�QD�4\�� ��k�E<��)i��2?ш8MX�ZN%�}$��4$�G}Z�� J�����A�3������w��t�`�ː3�n`(�
ƭJ{lEqf�JH.���C/����)�F����
Q�BU����:Nn.���6�6ދ���_�P4�����l���u�
s�����Xk�K�	���J��K[�|�|"o��#Z�yE����[B-O��e��U�P ; ��7�0�!�=<V��_2'p|���+<9���m����g�3V0���u���L��a�;.8���IX]a9E\�"�[��E�PG�e��ٻ���G�\*Qb�::*6q`~�'2�|حtY�?��1V��[���f�e��,ޘ��A�n܊8���T�&}}D�c�� �d-0+@�܎�7H����U��ꢸONLנ�ϋ@E܈4�\do�� >��U���ID��r�u��f���f?�A��T� �����W$�$����m��+R�(TST4!� �s0�\�!����;ӻ��:�u7�cw�N�Q�\cx@z��i��(�j�i�~�֙�HF.I���TuN5��t�*6��k�5>"�^J��)mnz�%j�ӎ�a28�d0]���c�l|��o�f�j�1���g�K8�!��T�$c��4z�. A�����I97���k�R����hK͘Uhk�U�!�|�����_U��"�-��V�l靎�?��[}E+�C�xekn��Zܺñ�h�i�ŎhaL���bˍH�w���gK�?ʋ!O�{cx�(��0�}�2��[Tb����.�D�\r\�t��Ab^6�K��h<#x��A��:�δ+��ZK�{Et����Q�]�Hj3��q\ ��2:7.&	0r���c�ޮ����3�%w����Ҏ�X@���a��Ց��eY��E+���!ŗh�;ë��ż�/�����`KZ����4�"M�a�nx�%�E�9٩�l
Ȓ��֡�)�8ث;�z(�x�jBw�ʉ��R�D�n=ɉxxE�4�8�]B;*BiSP�-!�EM�8?�]���${-,�%��&'$G��z3W�VDD	���I�u.�j��w.�/�|�8��n:o`����VMY����@ޑ9�RWx�y`u\�`������ �/���ó�~��p�"ذ�l≶�ڭM�$m����T�S��� Q��j�TB��+���:��V#�3"�;���G�jp"������'�D��~�4����m����:x%�y�!ʡ�ʨH�"�(8@l	;.��O����'�rX�H��	je ����!�Ԩ�]~�Kޛ~�l�E��\��)]&�Z�F����6:T�-"��X�
��_չMB�G�����hC�bq9�
��R��۞D<��6//�B���]bp�gj�5�N$x���]k.�ʰ�L�4>M�iLC���qP��@H8j��'v��ܶ]�#�������T�0�0:�y2��� A��a���Q���K{�g�b���ݝ�3�=����l�W��Lc5���`�Rھb���$t��L	!���,���Oɹ=~)l�OTԇT08�沭ԍ|�C�=EpQ�J�1��+Fdy�0D���a����?�YS�".�T��i,T0����������T	t���S!�[�'4�"K[��\�����3@ظU%��J�!.k���6��xR�[��ϝjIϙ��ɽ�&��|�WL9����'*�.EE���䧶��"��!-R-��#�*�uzE����:go��x�����@��V>�����/�b����q;���*�J
��O �,�<A�>���-K�rw�O���1����;^�ώ��M��:��������"����FU[q��!�1�]Ū�V���63>r�&���O�[�*H�b�����i���^�Y!�u��v(�/X9�=���؈�̘�Z�L��.��Զ#�H���A���E���oڴ���	{���(�5��_�o��TX��:γ5Ye��[拾	a����L'�9oq] c
L���:KU��Y�}Q<����z`�͂���Ͳ�M�PU�C	����@[�Q�P�z������g�Oih�mDC�ސI�u��Ǧ��6�|���W����(�����q/<M��u7��[��Om���]z#��/���x 68�0(=Db+l�K��K��p�scQ���Ɛl���Ty���K�4�͔�7������q�}�'�5th��X%�\ږ��,ى̶����0�ż�%�1S���z��ӡ�a�N��/�B��mm�Ƨ g
:��gfd_%�����;�����tg���z j����i��Z5�g66̨�<�-��'���Q{����4r�;��4rM�0,Gs�.�:F6��Jz %�_$�	�7&��S�a���DX���2�ZR��O���T�� @��sQ��`�	JE2����mF���_�E$�����0Nx�Z���@ۺS^��ÎRCb��9�����w̝i�H0&l3� }M��Z�\�]/��x�MA2��9��@ �=���v���ISl�9΃)��m�;��5~gU ���ci�����2���=�?!��s����`�.*�x�zn�燋��1��Xx�^���yM�>B�,�O(v<���� ���FJ��,/6v� r�����r�kE��!ϩ��%;��;n��_6f����ޖ��Nѣm}ZA�-�X(Q<�qE.�j�I�F��J�
	��ٴ���D79i�̹����n�1��M��&c&�O���T	�8A����t��A���ȔC
�O�Eet� O-���{s��Nn���ݼ*�t�M��B�h�?:t��� Ř�e�e���b_�?��SO��<٦9G�2_���ř��\�ɞ^6%���\���e�g���'��՚�N�f-��T��RôS��y�����6H�?q�e��h� u7� D !����Y�dY|����|���p6��g�sJ���ѧ8.PV��w	�M�{t���R읣f�,��C�iW����-~m}�kӧR��غ�{) sh�?
yt,��B"\�������h/3a��4��>�a���]��}�D���@X'%/~o6�i8�$Pd��K2�7�x
^=���O8��"t/�c,o��f�W��Ac�@:Z��d51�]�ʹ�f������2r�d��O���ט}X�]B���m��Z���5^L;��a�F��?7�05�#Tvt^0>S"�L�nHQ��)�t��B �j:�WR8\�b������1�E�����2]�*g�/�P�x�����늄��B��R��ƤVeU�Q	\����?m�w�K������
+��>��i�d��_n��6�s��x��j9����̒�v��ʯ���gt<�lR��l�m���Q�&UR�r��w_nOU%�l��o�z]D��Q��8?QW���F�
7���ա&���1��
��p�?ŋM{D0*�cH3�b�
 ��=u�y�Z���+p��̙O� � �^��LڇT몙�";�j �E�CW!U�l� Ӹe�$m�����X]7Z;���:�q�:ѝ�"5�qwC�<Q4j��x�a�ڮuq���p@�f4?1%�8����m�@Ň>/�j�{�c�OS�C�Ug����73�����a|���6_�/T�3�=��- ��5�IO�}���a~�Nf�>}�0|z~A�*$�jB;ԍU���|�T� ~��\d p���`P���EVM��`~h�(�C��o���Di�{�����YZ�zUM3ecsy�����eO��L���Q�Q����Q����w����2���X�>(6SMFF��[�u!Q�
p�z�O�\>�D}�>�����(S�Bi�r'��f��?-4d�	��pc��K'�������:m( �
��������Y���)!�a��S�;�ɕ�����˞Ns����� Z޿�vkp$0H�T�䦫���y
�/�����=�����w�\4�h�;h�Ԗv G�8��a�rޘ*|����L	���5�k�֘ss��������?��
X� ��)�1$���4���96��W���v �®���+����Ja�ܭ�"���߉�2����UHX�ӘL�Ǖr����-��=���C�x�R}��t�R=�\w�z���#n]�@s,�P�B8�זc@���١��(lq�H��9.9q5c��n��+2Y��t�J)�c�\���b�X�q	:��h
1Lk&��"��1v@g:+{\<)�A�Rf��>��|m��U�0�`���6	\��X� FGl�G�ˣ7�g9�ytj @��k�G�7��.Q���S�p��7O�������Uc��QX�^q�N1���5Ih)<\�c���S&L��]�>P����C[�"'��A�;ӭf��Y�ZFS_��V��|}FÝ��(�eo���hVڧwm%����d�q��(�98	EbXΡ�@�1~��?�=`�\��	��幃��q��W�M?�$Fj�q>|\�Y�]���Q��.�Ҩ�ތ�����%��(�¼]�
��.���:f��A�a�&q�hV�q9�	(�C��5d{DF�IP���%�Սg�����Y��܍qV�/ɭ>f�{��|��s�(7\χ�G��
�Y5_UYAO�Ю1��1�-D�H���H��OԈ(
'��J3nR�̥Q��|O���|K���]	ؘ�Ő�9��Z�Y�ų�M��=���t�֐ ��c[�Xh��3�AO�Q���i��Ⱦ���[�"��d	ֺ�u��C�Gã^��r�-���%򕧄���[�^�X�(���k(�}x:�sz�5X��S�q�c��{TF�+������5�ю��m����%��}
!&�����>�$��b��G��̖����Z��,
X�ja���j>2�e?�p���+(&��|M�/d�f�XlxV64EB    fa00    2c10ض���W�(X���N��e�F��]=��B��~�E��C��'�b�5C�s�s�!0#�nŏu V4kV2ŷ( �� 
�{|�103�n %��q��'f{������OFf_�� �r�h���ڀ��9M^�z`��!��TՉc^{�- fC�?+��#�����L����K�C�i��]4eFey6ۦb�LL��<������odR��E�͒�].>�ozRz�
�1=��"���ƪI��!n�18����q� ��1�9����(��n_�Kc��Q���,�.�m��s|���H@ӋD �l�hJ��ky���/ގ��V)�����8�����$Bz��AeU~�5�k(f�8�Ȣ�k��h��j?NS�����_ﾝTz{0��W2�AA�t��ҷA�zV�u�#�S�7`����v���|�O6\�1D~N�r�K�l�ZXt�khb�ڔ�C-b&~�@w��w��_��Z�Ɋ��ӄP���-��m�"�-�^�g��7����`P���?fZ?|�-=%p�ބ�I������;s�=�+����ڧ�wKP���8��OWv؁��#�[�x�kN,���8���(� >��Ԫŵ��0J��ǹ��L��h~�y�R��a��0��N�5�KB���L��M�F��|���5�#|���f�s&��`�V�	�,�K�a{�'�9�?uӊ��K�ʘ��4G$"��=>���2��	��J"hՋY��O%~�%*?�l����ŀFT٣� �n���dU㗡�x��� �1�_�y�)!nU�$�FҪ= (���kp&�1R]�}p���xcy�]�yBʐ�/ɾ�y^cm�uQ�v��p��T=�
8���o߸�ѯF���ȶ*��Z��z�����Z��w,���S��lh��Xs@-�!	Y��H�-pHEױ\g�!���'�U�]�F�ESu�7����j3�>p��.B��V\R�Y��Ć!�T�Ă�M!��4s`��b��� ����ԫT)Vu������.�7J�Ě� �iw���`�b��&�2�
� B���9dݜ��Z�8`7��d,�N���vQ1�.�1H���E���� �bz��+}�Գ���G�8�V��A+�$�����w'B���D��l�w�qdF���؞�ۻ?��i�����1ʋl��?'����V,Q�S]�ir(��Q�JC+�|Y�^�T/�m�K.ѫ0���E5#�aS�K�Y��	?��ɘX�m=Ge�
��	
��� @�K+����.f��݉x|2�ۛ2j�c�'r�p�ۆI����h˪��W�1r��==x��y��į�$�I���'�֗����"��Ң��5&|�mk�J��˃�I=;4�$�E���w5q(�I�$��}|�J_��7�dI$�h'�р�M�e5�҄b�4!��o��|V�[J�^�\a��E���#w�va��������t�E�aV
7�_�u�"��X4�ϰ'�F��Ǿ#Lo�Ji����:6���+�D�M*�@릕�]	��"��h����0�F���!la�ӄI�V��+�+(����y<�>�]GG��s�BC��,ua�����,M�D�i��t����w;������V��}ȡ	���:�T9;�Ȅ�6"g�����6�<�����B�n��X����f�T�pA]���ɺ��*ђ��j?<�O �Ѻ���V��g�dH�ۅ7K�@���w.9hX��&LH}P@c�p��i��,w�{�7f��<���i�p.���m�L['�Í��` �@kml��{���2.��o_��V�7���k�Q] òk~��2Y\HPz�e{�]k9�E��-g�o�&�y'���H+�X��8���A���7x��x�Q��0$i���k/C=���;��C\�z���{�a�'Μ=�օ��&�[��� �-c�;�U�ŪM�����}ɧ!�|�`x`�]#|�g�P�:��	��N���R2!{�v�]��)j08���W͇W��xa?��̭Ru"¸�����vԣƼX�P,v��˝�����e$ǘT����0�&,��F6�Y=&�����*2V���P{s,.�;f��e]���
�Ȧ��M�
�e���r4�����	MfC�~H��6�0�Ux	�~oi)۴�g��2����p�M(�D�HyĘ|]UYU�ܺ���sل�6�F[1���I��)��J
3�S�J�����c"̒OO�A�"�.P�"D��(����Ō�ɤ�1����`����ؑ��Ao��CoUu�!�pn͚�޴��P*>��y�5a֫=|)L�'w�q��2���T8�=>��`mr����/� �~���E�n�Đ�����A��s���@#��^v3NO+v���W"��zHX�������U��R�)ޖ�\��
�&v���_ӿy��H�.Є��\mh�O)Ց�IKz��8:���Y�]V8�=��ew��(�g��۝r\�����9�/��^,�몞���[�����)UN�Kλ� ���o��;���EP�t��`��C����O,��ZiؕC89�d{��q����GUp{����D${]�8�\�bRX����fa�l'<E��\ůb�w���C?���M�>I+��'�hb�H��hu������׼ًk/|qO�����Q��b�<�o痝z�iQ��#����Ŏ9c�����i�����c�'��j��0��"a��*m�k�����|��v{k+0r�Ɉ?�Qԉ�IC�y,�u� +	�y`�H�W�=�a���N�~K�s��1V#��J�����?:�T��b5�=&�5�ci�Y*�7t9>[ë_]��s�i���3Z��/P��2���2O<`�g���}ϣP���{=�e原�ڠ&����H��Т˰�-$#M�ڑ];��C5PT]A4�$?s�͑��\�������m._�{��Hӥ�(A �l�c!}>�ܢ!�{�BG?xU҂;��ξ�I�2>�����:�#�s����7k��o�}L�g���7 �R�:�oˏ�l�<��c��)5��DE�U��|���:�dU��i�$��?5���ew��>�� ���\q�4;E�z!7,�Z9�{���=�\�5.i��b�>~�Mm4~�^� �t���RHE)�a:ܗI�aK�p�ٔ�`��6�H�z�*���P�+�Lf)q�GZY��X��6Z�oA���>�]��9�o"��w��
h��N��&�\���5����+I��ی��h���|�O�	Ğ}:�LN�҅����u��]:��kND�3W�k�	n�jN�z������q�#�����ɝ��U�5�����o��s�̂��^yL�_��Z��2�G�{�?��1�O�w����w��>�U=�:��睹���ſ}��n�ܲ"�%�wLAo�0�97��U������-����f{�2b4�H2ѝDZ����T�p뗹B	�}w�	�8�z熔�d@.��gZx_TC �+l D�Oq�R4�}�9L�e���	�u��ɛ\8�F-����k:!�
8GHWU;vo�.w^D|��~���4����KiJ~Z?T�l0%�E�K�}XI��kK)�*_�t�$�q���.�5G��J�@Rd����[2^��=$���Z�ӻ�t+j򼡤�˹�b�$J�7�9� ���M�2�����!�������)j3�bY[A-�5i�b�+��u�K��-i��E Z��~@���'��CyY%�݁�A���j�{]�"�=�[߉_/*2��sζ;�)�|�3�9N$�K�
@o������ P��2ǧ	�Q��+�&����a@ߤ��{C�FW-xp'9��=��3%t��j��Uz^�dP~2��qV�QX�s+��w�D�� u�n��>���,@rRסY���������<�L�W��T�lI0*�(ǆad���Ec�V���eM��
�Q�T^�>pnA'tR��nq��a|��~�,#���}��0\��x�#� 􅄄>먊�[��b�A��+2֏=/�!>����X<F�p����Y�vT�eX�i4/@�,.�Evw%c�N�P��Y��X�W��ރ!�yN@N�]��a�b�TM���;n����E��U���:'ke�����sm�c��X	q�ɵ�.y���u���h7vrz���<B=�~s�J�{���\���h����m2�Re�Xe���R�$��i���tt؁��V�Ӛ���a)㏨07��ĽH��b}x9��~��xE	���z�_ݰ������ݵIB��N
���P2��3�&������ZZ��hqк�K���KN���w�~����al�#}�&\����6��vͅ�'qS��+H��2dˆ�N�E $� ���w�3æ�޲8'+.C~��?E�A)��\\7n�/�y1��v�E�*��-��˯R���5���ⅇ�\�BSz�rؓ��k�ݽ��PEl��JkZ��H���{t/�ok���� W D׀�{����5:o��%(~�Z��Y>C��ZaM/-Z7���̠��,N�Ո�@煰v�|��HvW���h`���5?2fW]��K�;����'���x(1����Ҹa,"��Cɼ�E�BH��n�6�v��u��f����w����[��[�L8�bc8���V�c���:Pi'0 (�@ՙs�][�#h�;��g�A�ud�v�����M��v%�U�b9�wL�ـ����ě�2�F0#㾀���(Օ����y��2߁5�byz�7�-���}�n�wqi@�W�G#6!�N��C�$z������
�� �̨"_���́5��_�p�#,�s��q��6�+u�1��PD,E�pd���֗�d�֣�a挭��N!�����lZ��k����i��Q���V���j< ��jO�~ބ�aXi+ȟj	�:�K���AF}2��� �wWOp�v#��q,-*���`wtzwΩ��E�d���)M�2Zt,�EV?J����@f�V�j�,�Z=ZHcP����j+�ig��؇�\������O��W�~|��8�5m��0�2o��Q3B�t�|Y���3�QV^h�tʍrA�v�w^>���k��j&:��eS�C|�m�`��$�|�k�U�R����G�R@E4�I���n�7BKm�#��X�cP�qYO�]Z����IDG�!�_�� !���tJg>�5<w9�~�ss-�B^?�g�F�2Yd>�>=�����!�9*n�� ����v�Э���zM�t���s�f�[���&
�Yi ��;)�x�����G��t�l�BБ��U;�U'�6�;D��\�ڽ*J4��ٓ7U�d:cHW�8�z�N�󖋜�7��#~+z�r3���K�xБXN�&\�#��S�RmԞӑh��^�_�Y�ѐ���Q,�d�A����j�k�E�]��ej^�̚ѯV�)PR��΍H�4�� 1���v���ȕz-�oț���V��e%��^_���.�5�ɽf���ܛ���BY>M]�OH�{x��l3v��
1�̛����O�?/l����jR�NA�q�|�,e�v��y��ڐ���a����7V�=]�u�8�>�=A�T�]>��"j�L�q]���?Jn�~ށ?^U�����a��Q~�0D�}��Jā��Ĝ|�4��۝����&��B�j�{��y�A����;C�YtHF�s���������vm-��k�ͻ^[�8���&7� ʹ�H!ʟ�����k����ժv��0hJ��hհ�2�N�L{k��k�oԿ�c�*���EE�Q�5x��͔<�'&i�o����z��V�ڎ{�齬�A���.�����W�p�䋉�����Άފ��GW���?R=`@�TA9wҧ�Vh#A�r�憒K���4wV��N5����*�̪d��v?�~JZ�'����~L��?R�鎸� �::��Gq1�o��B{+I��>�;y���[)�����{�u��:�ӧ5��,aa��A��SZ8��l�m���%.h�&����sz�U�Đ��-�w���~�v�����޶�N-r��ʌ����	h�G�ZS^ԗĺ��,Qp���dj�.� ���L��>�d7?<���� χ�:�X�p����!F���������e�E�2s�ȏ�\e�_�a�E[�3��ݳ����)��o�b#�`�:>=P����z(gr�a���X�9��"P��ˌYwS�o�ĺ��Pm�9]�7��nkC���|Ι����  s�$װ�������17ю�������l�62�Ck�A��r�,0��p��_���b��IF��z��?ƒ � �a���]6�[J��EJ���.����~3����$����M��5��uF�Ǚ���Z���7�3o"ߢ�k�U���������J���v�x��ꈳ�P��T��������K�@����Ç�T9�e���꾀|�5�pG�����CS0)�I�I���f!��b�	N�BJCnn��WZ"6wǏ��xyDyk���|>�������lO���Hl�
�m�m�!��l hht����VV.�9�u�����Q7��3v���	��~��-�w��
��O>�;>`�8�4�3@�C�֏@�w�G�U�-�b������2ey�(A±XBb7��+ ��姙N<S�e=�)Wӡ�y�7@��nݏ�4����(�
�k^V]|�~�:`xm�'y���k��=����^����TnfZχ�jA�Af:�|����X>`�$�c0x0�@�ޢ���x=<�� n�h�U�@U #����l�D!�܈@'i�v�K"�g����u���4ܝW��S��|�Z+M~�Yi�d�`?����g�p)���b_�f���Nв}X�ٱ<��.x�U���&�1�l��	[k�%,���nSEA�����>���/�6 ��SG���90W�ТU!��,Ɓ���q��%�'V����F��t=t��M�p�"�N���V�fLn��P��3��H�^'��T�E��������jK׫��Tх{G��b�7�'G�P�����q�y���	� �сX-��bb�2[&�Ji�S��kN��:�[�s�ۄ.��OB�2��hңdU���4���Wȿϫ�had�р먇��C�l�N�Q�+1%��Y�
\mڠÞ+� ����G����d뜣Rz�sfh�K��w�N�,�1��M�Kj� �+�w�..	8�zL���!��b�6�=$��8�e��m����@YX,���ݎ$e��g,�\$�s��{�w�E5�����p ��c,c�0[�K�	~���x�hͫ&�f���J���Wb��!�K2�8&L��F�,�)G��H��<K�+�G�I����0�Q�Wb������VSk�W�9�|���۰���G�z9']��ȍ�ή޶�)�Ep4+�PB��H ���t����g�g��	z�ȼv�w�⩭3��N0�(-5��Ɍ�������}m�}�v"s
�����D��Ă󞏼[��(Jٮ����6�OH�`���w=I�#T�ڗ�Z]�b����ϾLFK��W]�29�^{6g0�:.���4�lyLI~|�����?�h�.V}A���d́����9pW�Yc����ր��=��pY��˵�M�)Fu���4�h���ݣ�X$����������.��4�ȣ�F�z�9_������o>���) ���E�,κu� ����'���*8XruT1���E"6�:Mm����%6�F�9����5c~��7V#0�'��x��W)�[q�H|��d҄8*��k��&q�?PU)i}�����#��shd�q��iG;RH�'2D�lQy���Cʀ߸}|����ڱ��Ȅ�!��|i��u&�;e[���(�[8K'q��$)��)i�����*��A����g���c:�,|V	�O��U�a��_��5���r��������ٴ�|FJ8ݒ��s���o��� ���ӯ�����>l;*��!9��W�e��I؃�|Te'�����`L6��%	���B�J��F��Y8˵I�tw��ث���d�ѧ�"ۊ�7�^k��I�d�(�o�x	0��:N���ㆨ_��T��`?� �Dw/c������v�K��Cڐ�:u���JǮ�jݷr>�ӹ�&y�08��k���t
�b�ͧ��T�TqF��Ğ'gj>p��[�ԗ6�`�6��}�t<T,s5h!ܺ��w�-Q=?�C�FVDLd�x�m�686��I ��f�*��J��/s�@9�X��.�.��a��ݩ�\�UY-Q<�G޿ �T=�|3�n��(;��Q�p�:pERfRL�{�������p�f��k���ch��׭���S�~C]H�y�$���gW?7�E>����3�:�_�]��M��1{JU��m�Ȝ�{~�0�g��"�xZ"���T��Ȼﳔc�zY��)�jeX�۾9��UZ�Αx-�=��:ʭi>3�oĖ�Kl@y�-�C��`7�9���=����\���҃}l��/��i갈�AGb��2?ѽU&Gȝ���%�ѳ�ѝ���+���Uvቓ.��W��U����Q�Y[��Mn�PT9Df"���V"dK�)^�W��TBRR�j���|%�kC}�X��D�]�������]�L0A82��u|��Se�V��[�:T��9sȘ��~�
������Eڐ���{p��읰#A�]>�;�/p�<��рGg�MK��(>��w$Υ�^[��\����H���Q����·E���J�����2L���w�P���;GMLLr8*X�b��?��|Tu{"�s���Yn��w����7���J_ޮ<@�r�������o�ȡ;��8��ߑaك�.���k(��[��s�';��&4�+;�u�M<��I��o�j���u�I��2��E*�_9�v!� ��p{a��R�2� �ykF[��p��ǣ���\9��ܺl3q�po�܇-�Hzşې�V��nro��Soßą���Uְ�v^�O�T�J68��Թ�q;���h0��dZ�8�tF�E��[O
1�1���M.�V���FA"��J����ST�4U\2�B�CC�w��ˌ����rh�.{^�G6�w�j�i�]����(lSOҾ�`ֹ{����B�^eҐ��6����Y����E_w�Y2�sZ��86�M�`��U��2���	�bW�&o��ix*��"�pO	���.Eɫ�D��)Y�������9�M�܏5�B�@j��Ӏ �>��oΔ9T m��Q�;���9�x�*c ��&Љ�����E�瞮�9gD4ظab�f�1�xX<Zb��>��x�:����N���ѕ̗�pnX�)�!=x��	cC���aP�>.t<�8ov������x����⡒1B�O8n��~�����xƦ�;/*��7F4�Y{��X�@vv�'eM�\u��������L�Pԥ�;m�Xb4�gmZ�\S��[[x��6cK�?@�-�t07Xw9���@��6'�X���3�ۙ��;^)3�����ZF�4���C�6�X������W�c�ȡn��fw�@f����:�=+ą]&<]�����C�<K�ߥ~	�W,�i��:��q�9a��5��q+˽��7���s���K�`p�Q�Fe�Mo��c b��Q��� m�VfrK7l��^�yM��ú�[�!��%�o9�m+�'�l�+��<�8ܠ�z�F��AZ �ڔwl)C��Q�O�L�ܓ��')�~u�ݿ��Mð��l 	��!��>mh,>)�	��Gf�Ǒ�7xS?�X��:pJ�fI��&R�*�S`w=��r�Ł�f���2�rh�c���R���A8V�r�h�۝��Hu�x?B:�:[<�D7p���t�|>I����
��뷅d����;d)e��ލ v���杻�F�H���_
�ۻ��N�Y��ZBi�#��+u�~�K���o4���-ܞ%�/h]�d@��[CX^�~ھp�����/ ��ɺ�6g�k�0�>k��U���`=\�_z�`ϰ�|Br���o� <�����Nc%�wO�!T)���Ɉ/_זPw&���`6: �䦮}�n�/����6�(4��K\Q�}�����|��� ��GW��DÃU�M#Ӂ�y��u�"��p0�`�#'0��֌��E����	$%�@�9�XE���4�P ���h��z;Y���E�o����O;��B���h��_m�ι9��A�$�%k�m��:�����d�6�6U��&_���Ą�Ϧ-������g�����8C���h��]�G���y��+�e���s۩�t(���Q�r���sc��h��B�Ʀ�Һ�QR/���y^��� �̨������-�!)� ���B~�G�t�l��8l�Z���	:q3^v2�@s�(�\��Q�%���Gs��ձM���}�
� �/w[��oG2��]|bN 0i�#iWI���}�y�J�`*�*�s��Y��j�4��q�L��l$qm��O-��hl|{�P\R�k���9��ޣ�Z��5�3W)A���[\�$?s�+f�$���b#q8f'�T�}W���׳�^n��u�(,�E���6����jᴞ��/��d��g����o~/��q�|��Y���]aZuE�r�!D����vwj�]�Zw�CV��ڒ���صt���'+>���I-��c_mO�Ez�t ց:o���2���U����bL�:�<Һw`�$Qmpq(��2�ڸ��N�r��5FwL���=_��Pp|tM"�OwM	 봹�|��i�n�R�m�);�=�+��Bd��@Y�n��w�WF������kR.˦l�m*���{8��0�2PJp���-~BG��TU�@S�ݫm�א�z����a�т#���_X�'������|4�R���p�N�g���C@��!�?s����/@SNX�YR��d��Q�M�1�U����9�a��G�@JB�%s�ͮ�$8��	�]�v<��닞O�A����%G�~��*����t���E��4�����M�,"�.'���~An�0$��$.�E�'��ʹ�͛�u 75�)H��U	?]�99��q��D�
R:����s< �v��@���A&�l��>	�\�;�Be����Ā��_V���H�i���O`�+��rX [���	��c�XlxV64EB    97b3    1980�ʌ���:w�����GX?Q�;���Z	�.�4�W��	�����i���Yw���&�*jA;t��R��OS��8lo�i��23i��3H�7�d��X����ˍ�'��/A:>�#��$rc
u�����/8�2d�t��	t9ҲS�K�K�ʎ2���S�����f>��3ӈ_^f��3���ӝY�����;X�Z�@��Z<�UU��R�&���L{�܊����|M�-ep��
�� �\�z�!����3	W���G�{6[hn����\~̴8LA=���L���K�e��Uͼ.��/?���O��M���p{���շ2i�& cWQ����M��ҏ�r�#	�`y���m>��ݦ���9RЅ�9�Ӗ���������:�4���֦���tn�7��W��x��#@���2y�����ӟ��?�4iof߀H�4������`�R�r�e�[�]Yg��mi~��K��D�?�&|r�C��u�G��OV���q6��V�< s
��-[Ĝ��9q2�Ƹ-@x�N|�V*�/��/�f�F=.|�ÏH3 �
�����Zz��$(�qf�ǹǯ�t��'���ck�Of+���
��}8���vח2��4j������B�����̬#�i,�ʢ�ܕ�(x �{��?��k�㛗�� Û-�SCx�k���b�<R�,�Ŋ�*��#+1qŀ%�ė`գ��-�fr&P�W�u��E�p���A�j�o���	>��,+$�O=��/"zP�r�.5:�)��Ww�{Z�f|μp�I
"�=���w�Q�n�v�)��!�˛��(�I����ڲ"�gZ�yc4"g��!8�`o�J�xO�X���V�?5�[Lli�ۖ�����&s��	l�FV���-}�2>��dY9x����}�����0^g;����J[�����*��㟠��YF�-�Z�න�b'��#��ӓ<2�A���f�e?��|���2~Ս)v�$Nυ �����Z�8��GB̿��%�ofq�{�*+;NPvYl&��x��ڗc�p���T�م\4����&���3�!J�e�f���.5/6hD���������x���Z��ʚ�
�'�$� ���zPX�T]ˑ��8�2�9�������J�(�ߟ&Xp�.�u\�P苜@��}k����A��m�Р,$��v��
h��-e�S�r�h�	)�L�_08�o>Ӭ�(3��$Ew�拽/��D�G�K�����Vr��$�_s���:�g���?5qǚi��S�!�z~R�*��=��ܤ_���������E9�]�ZT7�!1gy����=�[���6�|�U�O��1���|���f���{n�Cz��S"z���x����}ӓH���	!��Ow���i|O��f����������>�
�I��oԠA��C�J+�N��7��<��
;5:��F��B�j+�65�i�)?� ��cy�&�ϲ�U�XB�{�u��p���jN�3@
�L�E��q�{��
�ҭs0��c�kxxf�=F隘h_�1| �X@2����{(����b9�,J�.����?�.��H�5)\A�T�nS����Z�!����,g�r6l�M�_6��}Y�����E=m!̯���ð=y�WIun���&Pk���W�IA1{��~I�V��^�����^�֧�u�0r�,h�j/����8E\
d]aL�x�I�(��D������� ���D��7Z���g�+��"i���@P�bq̹�&˝l|�,�����r��av`[Y]�D�����gPm�q�¸��{��+�����)ܟ3����`=k�K}G�R�-ą�|�Z~,q�&ށ��W�G,���f�bSEt�=�w�'ʒС�"cC��{���L�5��
�2
v �$�\o��МH����*#2��!Rt��nh��d1� \�J3A�!^�X�2���8�Dܦ�_}��g�m�t�2h?�g����=^h�'�~e'�(��d��z7�ힹ��6�r! X嗊�~Il�F���YA[N�ꤑͯ��X�ǳ`�`BHĹLZ��}��tF����sR��G���KE�H�n�L<� Z��]?�q���綝g�oH�a�W���.L-�Jj����@z����3���D=��╥�u�Ԭ��Ș��X>|`�w��������u�ZH|�ؒ2�n)\sj�K���=�ˑ���z�"-��C�gU��p3Ȅ�ٰ�c\�c�����򠠟%%(�B���)�:�WHt�� �}hf�b.�qt�bl5撟�#�����e��ܗ��%TI�F�M�#V�Anʍ��1��f�@�W�
c�S{Y��O�t�l���}7Zo��(��������u5�V���^�5���;\(�m����V�wY�}�At6��������a�=��t��H�mrO(>%�]�<-"mۯ�N�XsI�A�hD��)D�����?-�S��p$�^zL��&̚�rğSޓ�����fW��Ed[��V"kC�ܯfW��F����79���.(��4���m�6�8��pe�|�&ïG�p}8?���U��x�1N.I���h���d��a
ƍe�-@/�2��`��ߗ�)�9���]@�@O4�y:1�UA�*NJ]�4�i:aKb�x�o8����sg�a���m���o�>�ғ�k�n����gE�3��(�Y)jMH�T�;�7�x�$�J4�("-�{?Ž��&t�f�]����A=�5+�u3�^�T�I֮�-vO٦�O3���{���nKo�)<A�6"�	bX��~\�O��?����b_ȑUrRǓ]>��'�AE\|$ �����­�զ9�\)��pM�G7d�T�_�Q��>(=B
�(|�}l�>�Wɪ�W���c��m�B��Y��ٲЀ�J/\��_�4Ch?�?]i�E��E&z�Z/��&6?m�F(p�ª@�>K�!\&၇=21�c�y0��������H�x�`dH(/��
�<!�c��RۏQ	C��K�Ɔ�;7��*�=*])��$V�y*dSm�)��N����-"l]X�E��?�PP�z 쒮s���IT������d�C�]n�`�t����_���A�oDǕbJ��1`ό�n��E+�E�s�����s>9��Ր���ř��M�-�ȧ��܍�r`�4a��݂����=!�H�;����+�	���돉r��N�q���s� l��E�L� _�N]�_��5߲���l�;�\,*>�Rɚ������a���ƙ�^�-���h�4x�_�\�6~�2���=�*��t�<�j����^~��c2����]1Y�c��x��D�ۭ[�NW0�vD�!���&�3}?$b�?_�iV��wm'�f��� �]�.G�� =�[�IO���+4t����XHJk��龯&Wl��>��K��q���W��
���zܼ��ʜ&�Z���w���v8ӻ�e�*�a�����y���w�\�_!V���W��F������]8�q7��y�n6K_�T�(z��zU[�b�X8n�ֿmM���7�COt4zfwC5��!DZ�)'=vc�����s�,�
�~y�$K G���tf/�o'��Z��੝������
`]��������o��tK~�$��Q�Oӳ�?�9ǌ:�l>��ظ��C��#���{9�>҉&	��8�4fTwXfb,�u��JLԀ��=���#����_�5� ���1�(<w����?�4rޢD�X�0%j���~r����DchL�,��ш�d�d`v��xl�S�{]����.�خc`1�mk�2��}GP0{c|Uk���sЌ!OK���5=J����\��yǎxp��J�K�b!^�H��h�v;:���([p�|.�nW�!�m��te�T��	P�aI�)`8|/1؁ܦ�4���6x�;������5Cy��m]��ŀ&�]el��ؾ�&�s��b�a�2t�w!"�� R�t�a�����̜��_��>��W#��Bx����H	�~���G��g8�^��"��ޢ�}���]lxT A�h��{�'\�:m\���p���j4��3�$���SMl��X�}P��ج�5�]6�5��k;$�1��U�/S`Rұ<��͘��%Q��&�M<�����q1a�K� �gwNn��֞���ڧ��JI�yM��r��z�C�7��wY��Se��/�[K��F���'�b�77ѯxR�!a�VC���?p���.���c�5������;�r�!��'ثv�Hw~�n�d���z�#9Y1[&%S:�K��o*_� �.[�{��\u�U0Pz���C�Hj5ӾӖ�x?�,�kjX��=�s�ڄ��<u�g\,�ۀuX���
�g�F�ë�)R�c�j�&��T;K$���Z�ʁJ���B���n���v��B��)�\�;ZI���dF�>EF.�T�~�b��D��Ɏy��Uǌ��c*E�M�.p��6�1�Cn�͕����9�r�����t�Z�o���V�C����v�B��0�Jtn���vڳ�r[/5�h�o�&y���-�ݟ'}�F-y\���(�DSr%ѭ��sV/�5z2�\������!�,��q��W�g�$�M��c�ʷ�k��V�_M�kI`�F�B���Ф �xv���4����բ�o9��m�^�	C|������̌CvK&npcDB���o�����*�'U>-赝�����f�MO�p�}��Ҁ�s��g�}2�k�1$��9���G%+v��m�
4��٨���͝%��2M�A1+�Zj�zyw�[���E;e�����Xg� ��?9�:`�E�s
�����EU�	pZ�v�F6�a����;9UTl���=o�T]��G����y�K�6`�X����ʾ����ȲmGBnη�7y�7u�����Q����Mf	�P��󪅎�b&���G�|�H��LK0;���Z�� *�h�Yв6f?iH�(3�%Y��rw��x����Cc���]����Km�s�xF��c]�>,$����E-����-y��@J�����q��0o�y5u0�X3�&pm�[��?��E����n��š���̬�\{�Kέ�ҽ�y#�)NV���������U�=,�a�@|��������Xm�n�%.q>�+�r�i����Ltc����gE�ğ�h�+�RR󹭼ώRe���� �[Ϻj �`m<\�d+x��4ȋ!eãi�i�Q��u�L�K��￳��:]���?]u��K�Ňb�U�:�'�� �󅲔�}��D�>\����਻�  �21��g�Jk�:��X�t]��b�6���3`|c`[ʩ��	��c�/�Ni���D(��3ʁ�*_�|-?,	ٵ��Cz��4�S�\�ۄ�q��P��Zq|%�az`�M?�춈-��K�2�Xy���/b�F��$\��x������%ME���$���/}G��aIf� kS<)��J,H�g?�d ��h��'F��q�_UD򭐅>���3d*3E� ������F(��{�0M>6X�v�u��E��aӣ~W��@����jK[��K7Ȭu�9���a{Z,;���{�1T�a�NQ)z�g��?N"K:e�M�&�Dh�x�g�KEž�j�W|;ؒ���&k]�Ԟ�>x�>7k�R�n�Yߗo�=��'�>�|3T4�nǖ�����F� �'�[%~�
�'p'�{����G
7�C>.>6
�6��m�N08�L3Et���)��k���K����?,�3�~4�&$%�����{�sB:�[
���8w�e��*$�3�2l�&����xz�ʖ:Sd�6�4�ҹ�'�c�<#O��H�<�U����Fr��\;�E�_^����-h{%G7�=2>��z����[���$�D6mѱ�Q _�찬����V%���6`��ĭ3�Ѵ�j:-����p�h2�ɂ�WR^��\�VdP���
1�J�Z
�l��J�*�VI6l�8h�*�r��W�xi�9��#�\$�$����3����Y?rz���
[W���+~��Ѱe_�o�V��ʖ���w����Yc� �=>��H�ƅڑp�Q���8���tʿ?��4�LĐ�cJ�9~Np�:Ũ�w��HMщ�;���(�{�'R�zZĞ'�A!�FC�Z�ި#�'IB!�lƌqb��J̌�����x!��@q{�"e8D�L>8A#��\|�<~}s��'u���G"�����F�˧2b���av�1��+6x�+[͢*H��#|z؍�ѧ�m��Ӵ�2�KE�� ��(X0 F3�}f�A���qa#����ٺh̦oK.����iE5�x!�`���к����
r2����]i��YA�ƺ�2�x�oOVja�-�v��,L|!�F�@>;���8��mj/H�E