XlxV64EB    b70e    1bd0p��B���@Wa�L��y�	��V�ӓE��d�x�s�iV��XR�	]�O���`��ˤkY���"�<�g�F>j+�b�����P,�c2�ʏ����}F�+�`Y���J����\ǆy�?��El�(_j�/�C-�I��ʈ�����Tg(}��d�{g�:�_�h&���Q|�+4��ψ6j�������}�L��>�05�&�[Iտq��@�;�┆���4$4�Wq�˧.�c$�>�C�*oE�P\*h����۝����p)fo�wF�y��8�Da,�F^e*��{��~�{�xfI?���vf\�].�j?�&uƶ?�gꎮ)]8B�N�c��ٸM.F����w�	�i�o-t�k�@<OlĻFD���E�n�O}4��Z��28E/:,��X��en��ZB3g���FB��C����l��b1Uͧn�̇�� ^�����]�7����TF�\� ���@�뷑���˖��!Y���@0	���iù������ڂLh��3������$�}��$�ch�u��?]�3s.z-����<������ ���uu���e*��%���2쥧��>�@k��
� �M�LZ��-��(�-H��8犛=�')q�
���(���8[N�QՆ=�gC$XL��� �@k� 	b2=B���Sǩ��rŇ��2����P:|���;��̌0��MY���~�0�F��9���m�<q����Cx��a��]���#�T ��y�K�6K�s����$��������u��H��[S��#Y��q�=y�h_�������9��K��M��6EvS	��"Ȟ�Fz.NW7DC~jζ�2��)V�X�p%��Z�̇)���U
���N�cg�єYiyYK���$K����S���#8LT������ȕ�^ߴg*�t�ӆ�9 �3��9߅�R���w0�����ds��{����Vܬ�nc3���R|����Qc�;C�$�������5������;k-#>2�+<c%�cLIo=/#����i��Y�a�Íj*e'i�0��ꓡN� �Rb���Ym��fy�vR?�B�2�%���&F6�m՚��l���`�?<s==��A*�����%~"V-u|3�٫yE�ڦ��YH���|��TFc��@V�����X��.ֱLet��N.�,�4{K��?���LH���\��ً�0����`Ϥ�kv%�Uǌ���{�6��--�����Kh&��҉@���S�=SW֬jԉ�e@�Tڍ)�v�ښ�v��~��,x����妢;0��e�Z�� ��]5��k��]X��J�ť�z�5R%��on�o-�%�%�ls
h�`o�=~���g����B�N���u�5k��f�1X��
-&�-g�����r�4��:H�|u/=훽��`���z|������	����B��3��rF}j/�Ԍ�%�zK�`�G�o��P�g֭-R�b��e�Ġk�̱�u�d�9�Me�l����ŵ������?C��z��=1?�Vwa6�*�*Y�F�,no�8׽f�Uo5ʞ���*~Fg�&T\�$TN�!o9S������1QC����>jť�{�%�bYݴ�C\�eh=Acޚ��{@v&Th�à�b��U.�����0F�Էt,vʂ΢����ߏc�������ݙ��V��l��Ҏ�ٸ�TW|�:�*���i��X�j$hn{��6�\̈́��'y(�x �%Ϯ���b��-9�8R ���C2�:�r��/�ozP�Ϛ`�����c,��0k�H��L-P�{V�}i�����P�����H/o(r�L����O =%��L�RΟ{N��%�h4_&��CcH.z&�ǙI9T�kze�x}�b#)4��)P�K ��Z�9�ٍX7Ql ��v+�"�O3�C8�@H�Q{�
k�Q4��}d��[15�#��)�U$��|�"�0,���$�� r��>9Q�3L�SY��qK�_F���c|<�	$�m4����fl�2�l��#E��ߺkk����1��ܖ}�����T?�8׮��������VZ�JB~��p5�w�`��Ž��25���ధ�E�Æ��>���}Qʺ�c�߿�Ia��̈́
~+�:�G<���^ju	~7��������&�j9���+_�����#D��N8��7$>gk��������S��a�ǦѪ��OC,^��e�����;�HFX�g�?���m�x��"�:�f[UH��\�X�d����÷��Z`,Vl'^����Z��xr!!HeE�6ƔM/�6�:]��@�L߶qk��V�W��cUB�R�����v�x}S�:=qA*���V��٢�;[�{yn�Ւ��-��C�0E���D�o�b����8�#���8�%@�(�P3��*�(l/Jɑ�61�X�#��J�Θ>k�]�]�$������.��
c����2��r��i+���'7YyV.Qs=�J�n�?��d�(R�V4�o�3r��`EG]���=2�}����<W��-)Bv��[��/o���e�	�5��3ӟ�p�I�uȄ�����j 9~i���a�7�E�Cq�����۩���˰�M��8�*��^��SH���"%�EQF^^D�����bY*���)��vL�P��� �b,�@�cpȘ���[Vo#��\m2y�-H,IV�%�1Vg@PQx�" 0�6"/�ח��m������0� v����0۷��1=�	ZߗG a��i��v�F�Ȳ#�*T~�kaP�J���AY:U8���iK�R��
|�*ʙA��&���̀o���!����NQ~a)���Ð���|�S���p�w.N9�W�)�8�Y�KW!'V)o�l��c��u�,t�^nж0>�eݜc����v�_�"�e�e�Q�6��_�.�tuӵKP�Z�ˎO�MA�����ܝ����@-�R����
ҙ���қ��s��UWT��Õ�~-Zg_��F#[��7�ê�qf	�P�X�cij9�4�~�7�J+_���*Q1"������b�L�99<P�������㌱�>:����R ��,4����Rb�#�����b�h�I�Q��|^%��,� �cԍɀۤ���8d	7�-6 I��[3�K��0ʱ\�{2�֜�aZ��=�~�p���i|��Q⁤�λ��	�}w�`Xz���VSu��M-�� ε�ӁMl�j�C6�Iٔ�<��h����=$Gcb-`�- p��!���:���_��TJFv���i�����<�y�@�v(}M/U��4���A��!^��RZ�#�؁ܬVn�;DA8no�&��֗k6���a*ᡖ3"�}W��K���+q���{���G�3�?-��6V��$	��*�/��h�����#^E8s �)�e��do+��A��%���F������<Z����I]#ۣT�%F�@ɞfbR�΃ǕCھa.�q�L�}
E�8�ٗ��5��h��߽ƿ ܪ�� k3����Sk0��h��ZѢ<ǲ��X�;xzv�<s��y�]̪�{��i�;V� Ц�Y�R.�_zV�b���u�W�ͣ��U����,��"�(0��y妄��<(q�h����#�"-8�Y';��O��)u0���PDp��ձ:���Mf ����[��U�~�"(��[��k��q�ǘVݓN�* $V+C��H�'``��#	8F��^�we�e	^yaH�QD9p�$::�����X��E޶0SB"�9K��RF�q��N{.2��z���ʋt���˭��Oy�	;�ׇ=�̦�U�����*��Rܜ��v�T>�+i�)D����s��it����R�Cdl�83�I��.8�Lt��H�l+s��e��CGw�хv��Rr��7$cͥl��Xt����|Y�/f��%�L�4�H3L�d.=IH��$�����=c���x�Hq�t/(��!Kyfd-�4ޟ5sNS��?��	�i��OO�D��$?tb^�c.'������O�B�]�������`�����׶���9M3@�)��Pt�Pt�:Tw}��RVj��lf����J��ᅭZ&��Zذ�-�@����.ބebv↶+�S�x��;�V��&m�z���-����A�K���N�`匳�Oji�^�o����p��@��Q<0!f��*T���I��� �!��Ѽ��9�n�z7�/ۢ�&�|��S��Gi;�K	��~�MVde1Ј��E�Qw�J易j����Τ��E��%�0Y�>���q\c��J9���D��CMtH� R��KN��P�J=d�r�JT��ox�~vm%aߌΆ��.��ќ&7_N�Ck���+/>�ֳ�El��8��f�+����B�JWl� ���Lb��L��VWE�ᦜ��^FI���޻i��8�'�ª��x��d�٩�)5� �fe�v0o/<�0�M����u?���C����4�,~e����6��A1��C1{�ۊ@�fxo��.�|��fr�����Y��|��&{w��h�џ?�������}�ΔCr��=<#��n�X��E`(;Ɉ~�m�c���*�J�:`iU�t�a�S�B~fqu���)S�Mo��&����������ӄ��a�z������t�x�bJ��46�r\{h�\U��Py1���:�r:S3���Uu�4ޒ/��^�?��Y�_>뗪�0��Mz�P-s+�U> � ��r]�	� �{�;H�O��dGK�Ǽw�i���c[d#�]�T���#N��
8����LqK�p�Z��;�짋bD4�N{Q��+Ū�p<�C|s)���X���W��XT���ʵa����DL],'�N`hb�i�^����V����SjJ�9�E�Ɍ��N�	�,fP�ˏ�-VJI4�����ʮ��i
�#�my�.6�����Xm�b����iҼ���ң�p8�,�:��m�����.������9%<�eb^���L��ع��	�"���$��9p�<N1,����4!7���8�e"�5IY6�GL0CԻ��:.�+�U�Z&��\u	u����57W��ѻ��_@7�� �XRҪ�txF�xFp�����_�k�Ãr�m��:��oJ�&0z�,]�[�X�-�E�n]Cȧ��4�[b����z׊= �ay	�j-�/6�J�/�n� �>�/�2�X��(��(pί,��)§Թ�ӕtx�L@�+Y�&��]�l:߇O\���q�����^\d1jX���5ǡIVm7�ҫk�1�_'��\�UR�R�X��λ�m�(k}�%L�BQ���Y���Y�T#h�t����ʖ�:(��<����M�D������2�;�>l�0��Fh�m�B<O�o�&`��n��TZ�E�Õ]K_�Aۢ 1r���:�^REL�T��וY�8��� �~��ؚM��/�Ҩ� ��؆��
��'.5��i��|��3�n_5!�F�p�؊8�%���HKǉ��ۂ�WQ8I ��Z葞aO�,:���j� ��Wt��5�;`I� ���	���.�����a��پ�G���(;[Rw>��Y5C��+cpF#�&Α�I~I!P_y)���A��M�$���4�[�tp�?���(�D�QD6)�.��&��sm% 
kC:��iS�� Γp��O�#qY=]����h���I��r�d?�w>u]Tjj�f�E�0%	H�)�gp�*_�9e�om�`�)癫G#%�o�i5C mC�����u��пw�J��ٶ}�@������qR�1^��H=�����#�!�aV� eD�x� ��[c��C�/�)����Fy#�G��B����4�y�t�(�{nؔ����%nNڸ���BL�]��z��:Bі�j-��vi3��n��:;j?vU7t��Dn{
���{&6��:�@~�t!��و�/02�pYem�ʀuWw���jbӰk�b ��V��X�ЎVQ��SI@/@*��#��nt��ڡ������$�0����E�[��o�~Q�r�?��d�G�=|�Px�K/`zB�����;ws۟+t�K�3�Rj���ɸ�?�bO���JA�~n���̼��N�5�S��N�<�Pq7?���Q��WY[�L�;-��#*+����?v0]�}	�]�8��ܜ̬��y��<؜�JIz��ʁKPc=7�����8m7z�"�N�6]3�x�q :�_��Fi�S�ؓM�����g���:^�d�����,�z�?�Y^��^���X�o1��>��Q�av_g,0��Vo�Kq�H��?�����-���(�p�u��~,G��i��� ���:�q�4�|�o��r�M��|i`���փ�������bl�M�xź5�	�3 �k�M��������
�)��=q�C��74K�r&�n��M���!D�����|�Mv�'8l:�D�gFn/-��r��Ny�����	��\?�/v`��|,D��Cjs�GA###�z%�HT�1?;�}L�lp�-'�- ���+����͸v�qS��.�Ğa_U�+Ԅ����E^�F�:�� J�9 ��]��g8U]Y	=?U�/���:���:�x�
_c�<�ƿ���_4�Tӯ��&�g�Y&P#��$�"��u��B�x�]�_�Ul��&���r�k��S��M�q��|�¡&�%�5=���D�w�k�y�dPz� � 	��0k�E^<��-�f��ݨ��6�lQ��萔�͝�s�Ia�u��l���r&��8bΒުu��WeM\Mok{�R�i�U؟da��	��,9��,z��o�����jO��m���i�z����p���qO���3����������Bc2H��dԎw�a�;@Um���*��GX;?Ŋ�'WK�܊j�*p���,/����f�����(̟�	j����es����N�3hL��[c�ŭ���Cc� ��!yR���=4�;\'����_�%F~�����K8g-��ߏK��-FUD�4��/