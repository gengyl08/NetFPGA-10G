XlxV64EB    6e3e    1680=&a�ycVM��|�,�c�;��6���^m+��!��?j�;e�~)	U�OB�k���n�n$^�
��:ry�0�/���=�x�� �z�J(�L02텝Z��? �E����(��/wd������[�n�#�E��L�J�[[Yp�1I�k�㲳�62���4��cd�z�s�D�,{��j��_l�W�f3d������X�@KC�c�!)}w�z$�Pbjc1�(����1rxt�Cnelbg�\$���CG�;pykꪣQ�"�~����,
oE���)�;��d�ٖ�v|;f���V�C>��y痲/��I�voEE9���	н�0�@�mh�g����+O]sn�m!j��3���}#��B�i�ɋ ������:�J�Ы�Y�z�	R���ʓ�ɖ�)}
�-
_� 0�n������/��,��,����zڗߺ���q���7I�ӆ�#�g4{�b��B�vU��@�}+˥�O����MS?�_��� ���n&s��Y�:IbN����d��'���
_�[����D�j�����p�����trq��}����P��=�G��&A/�4��Yr����q� i��%@9�9�����vNQO�d9��a���fg4'{�<�p��ӱ�R4v=�wt���0n�'/��盗FV/�K����2�2�9��<���»D�����J�_B��'�R���4O�g��
w�0,J�ǽ�ʜʶ�1
����:L �I���}�r��a�ƥ�g�1��k�&��.m��"�o�~+���v6H f�YDwT���-
&CX���Q`^�J�:7Xjy�3�I��LK��SO�(����.���'�>��� �:������/9�\��2��-O��H�m��������:��;*mJ�e��¨�݈S��Ûv��_߆N����kزnj������L�~��jL�cI�3��@����m�R��Ӑ�~f1���Fε;VO�/$q��뫝����E��"8(yOr�FIaF���_����y�V:�>�� ?�,=����ߧ�F ]�7�N}��U�������_�Y��Ĩ�ro������G�]_@��:�N��~f ����=^7UU%�j敒<x��b}�6	Q���J;��`���O�z�2g?�(D��ՙ�������"�r���Ǹ:�Z���u5�l���wOM~�òL��Z�T��U��M��W��huN�xkk�I�P,�Hͳ�NG��ʪ��총ˑZ���A$�%���Ҁ��U`���������Tm��I�A��U� =_l�;��*͈�9�2}ؾ�н%iX���d%sP3��X���7r�D�D�ǅDIUq�����M2\���Y	qZ4����5}ץ���ǭ��n�k���@����y�N2��Mj�?�&�*/�}#��s*t�&���a,1�3m�<�M 5�;E��A'�8tZDk�h��&&�d�zad�J���!�s�y�G�9^Ȯ�~�A�^�^%Z���A̫`�Px���:<(N ����%+�޵D�|�����\e��Lzcy(��S�QA7u��Q ��l�2�i�|1�ÏD괹u&B	g�3�q���f䯏�
T~�m�uѾ�o���㒞�脍��
0�F:ٍ�-j9��j����i��E��n��VS�>`�6����$v�b�-\ٔ��2h�����[����^U�("���K�1���`$���WYdL�������EIm��O�k�p1��77��d(4M�*�5a�N"(�Z#���%�}W�$|ۙs֪t��d�9��ԟ��GWC�߅��e�kT�%�	�!�J8o
��z�>i6 c�	p�En-���B%�[��3�#v���p{�	�F;R�%��r>F�u���~�sw94)�)��q極-�T�k�F(�%"-T���P=6�В����M�O�C7��	O�V�*-�8k���Y�ґ8T��Ume�UCq�B9������zܒ��p/+2��GӞ�OR�IΏ͵,�"c�)0���I��Ek��ai�߳�wT��>V��7F[b����o�x?��%�~T�aY�/T�aS,{ �F._���Ū�)^`Exj;�ok͞�Z���H����5dy:�H��9��#��
.�<� �J��NءR}�)�n��b�,~�����͋��EZ��>�*P��GU�#k�S�eC�/�#��zzJ���m�$e�d?����ӗ��-Қ4Ͷ��n�&��E����2q��>"b����k?��q�:4�
6o�����us5�7F�A�Q��e�}|'�����⧯� AG ����X8)ݕ�ʯ��F��\O&�4[��3䩔Z��t.g߮��}&TIZ���S	���sqY���8�a�?�����7h��'�W>:�tG�xG�d�6ll;ūK� L��f>�|I��K�,L�.�WZ�إ6m����O��j]	&(�a����
	�%cRp-���2�RW�ٵ�XN�7v���|����	��X��%� ����BԶ�|�j����`��e�Şv̏6'�rq"�����B���E/7��?֗�'!�6	�z�� ����H7V��l׶�Fs��)�Y��HDF�оE�u(s7�V�����oീ3�B-�6d��Vp��'��,���V)ǴE�LDg�1{_��>e啀ӳ̢e� ���`1���+�G�NZY����B����Ԩ����|�'E�y!�l��o��'�E��xN�D��{��=��?P�����Age�$ص���L`��-�v�H�pA��ـ:�p��V^�����b��E`�4����v���~���!ɕ�T���!_�"CIp����΃qm��Μ�Ɖ�Ey�b-�Ɇp�F���@�`����ʎ$�Q���C�]R�]�_:��%q�K)7ɬ)�~[���MCk�H9]*�V�(���#����{a�����~]m��#�I���H��>Z�f��K��֐k%��"a��#v�G#h�І����7u��}`����'�����n6@?�!�d��6����L�?�G=q?��P9-Z	���\�=�Xgg��aT�ʠ�<"�͒d��a2{�~�~��ien��t/�*�wn��6�q���XPi>8��=�Y>���g�>l���+ٳ�
̓���A*��%��y�aZ�5�(�F��ߡ�z�6�Q\Y��F���hӉ ꠩[������X���:��@3VKi�h_FA�NvY0�,�'. �9M��u7�O�`2S�Ҷl������{_%Aΰ6	�[;��1Q�Y#�<���2��&�d��K"��e(��f�O$`����� �sw�9��E��sc7��?a?Z)mb�8,�r���Q4�w���i=4�g�������b�����&J|���J�e�V�b���[�-j"�a_�Htg?ԋk؜�[@�Dr��D�Z�x���{�!g㮋�C�������xrd\�dk���b��J���~k�=��W(ƺ�=�I7C�%�k�.�{v���ϭ_l�:�V�A!r�K�Z�r�}�@���R�D*Q3�����[��+Y`&�V{�x|��z�� ��շe��<��p���bwe��
�%v�B��V��N�n`�-[��n3�6R��Yu�`H�j�6n�@<��V��-�ٗ���i�#�V;���� ��������PC&@�:ԗ8��ĐY(]�E�'Y���~<�J~Rzn�/G��4��p���h���fU��/_�#�A�'f�QP����*�Q/��!���@�W�����i�木k��&����.�P���96�~F|p�xTQ�*��2�h�!i�����۟�!�ac}�rV�?	����b���6�scYJ�Z4T'k�ɺ'C��=����$�C`��f,X��Î�4��-��ޏ�KG� �l��֢b�����~x�E����1���K�D�m��]wq�3G�Y�I=6�Ú�	~��K��O�/��5C
��%�Dv��_l���N�ưx� د>�v<혥Ć�����sWx^{�t�c����;褍�l�����ˢK�FB��4�{��o^j���G��]&�l�P5hT�y�Gd_O���]|�mVח�G�� ���Z�ǰ�����q�+@2�T���`d��/p����b����>6j�����)��E�Lw�Ϋma	c�;���0�	7W0\5`���yĒW�s�h^uf{���>��tXZ�;F:�3�Sy�W��j�ÂJ�G5z��E>�as��7�l���� ��œQ��˫���J	��d�#\u]�2S��޹��޴)�@�*Ʊw��dY��D#&ހ,6J	.B��7^�2��ν���:��˭�������:i܋\A��kj�A��{��Jx�T � ��؛C� �����TAm��J9[���r��,��W�t�U��J�)���
��	�._:�('���HϷgu���[�^�,(\tr�w�8�!���:�����P�bCe��5�~�w��1��R�n�$'����*?#K��8=�EJ���5��
R�|���2����ծ�-j'�� ˑ�`t��?F�����,H4$�~���	U�Fy���Na�"���Ǽ���O���~��:,ȟ���p�~��G��L���oTqe��Mp��T�_�fn7�h��݃6xk�.̓�!��ћ����} ~�3M�:��fw�ż�7.��ȕN%21���J��� 5K2u?�^/�z(V�{���/�6¦�L`�.̒-y�<.)�U�`h5N{�Tݮs��|@�K����X���C�hZ��qif��
�V6��`��o�ޢmw��=�� ��X���j�����=#ʪCp4g��m����;+����T�2I�:V_�gG������1tg���Kڕa��:��Û��$��*����t�j�qP��B���9Bt��D,%F$;�TO<VG=
��k��x�4����#hcO���c؉{���0�e���������]�~��oQӐ@��Пu&���@'��R]/�1	�4�Gc�1}q��1Ĭ�h�V� ��㩟{�OEZJ�=�ͣOS�ݪ^?���a���Zk9�d�E t�]�բCQH����E=R�H�YQ`XX�Lc)+�<�_?�uA�\��@GM�p���4;!:�i�+���:��� ��WT���btvL�� �{�1^�Gs�ԟ�z�GN��Y�^�b`e	�"�����^���򨟿��t!���!h��0�z�l�L[$R�#x��A �qT�/ P��/ӏ�q��v<�nZ�8�2��cwbjH4���b��NQ8��K@�ߗ���#�e�6��Ɇ���Cs.�1{����F��� ���f$�f��X�`�!��&���$.si&k�:Q��Z4.]��_J�F�:���Kj*�tX�q�hn�M���`3O���E���b�Z{dU���B7[&~B�W�P20��T�����B&k�j]���}m��1�\���#��*���Аs�J1k�-d��
���I.�ϟ�����O���9%�I( �X/�0�*0{�[Mf����h��|l��G�9��ْ�G�W�@#u��'l��z^�O���sXƻ�Bh����W��J�	�RvG�y���[[ ���m�ѳ�`����o�U���Y�aj�k$e�{3�@e��<��O�K�S