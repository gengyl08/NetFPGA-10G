XlxV64EB    19b0     9b0����n��ka�� �� Ԝ˜��PG__F�^�-�<�Y�O=j~�a�PuJCS!����N�[�����%*3%����}V$-C?�2��e� �K���WCO�o�$k��$Eh�E�߫�t!2	l^��2���o�#5LL^Z���L�(fT��9�K�{���x*����/6��*�BM���ІT�l�1����s��d6�}�����|l�Mw%��=���U�����W6}����d�N$UD��Wtu��sLSo��� �����{�*��)Q���Z������=H��p
lE�ɯ�W�w�v�@[� ���|G��v�fj���ąw���.�ܞ}o�a��A��}A��#T|7taQ1$�|ͨ����o�Q<��e�?�<i�K�M������@�eF�#`g�' ���Ѡ��e�J��%B|�e�hqՒ�(��}�|��%����z|v�vWch �[�w����k~��a+2d�0��q>�_d��b�q���e4/jbl(A���w�9�N���9��[~cU�& +���3��3��ڣ����nrLpjp�ė9����4�����w��On�@rC�\}��i�L�Y����h������<�v�c8BA�%�@#xC�����&���B�"9��
�q3:��s��Ę�\�o�i�.����h����zMm�/�0�����(���p��Z2�A/i� �C���C�ؿ�j.ѓG�Q�T�گL�X�#Q4sDW�FL��r��9"�nj�	%����n�7 ��X͍���s����ZӃQzX\�Ɉ��#s��\y��f�<��aW��ogɱ���7�����cwMoo_2�f9�a<d$"x3����k_�@�E�F�����t��I>-��{��!w]'�Λ(��9�?���4��F�9���쥃D��n*�W:��Tr��	:m�����b�<�!g0w�S��=ˢS�b���bD�ӭs/Sf-��
[0�b�ژ��0-;	�/�m72��P �$F���������z��H� <I�����Xz9�|C8x�P����;�XãY�}��uK�)wJ��BrP{
�(̒�T����C��jQ�|�����u஧u5��J^p�,���p�����`/d�F< ����^�[�$�]�lQ/4�܋N�>S�h�xuڒ\�^��gU.
`l8��A�m��<�t��c�K�¥��8l{��>��ϥ�,뢇q�/I�=4��w���pT��٩i�/�֥v`���j+�!thO�a�l��V\\��@��K��M�I���%m�qS���u9W�nh�Z���'��.�uP�|�j���j��5��/��OԠ$}��ߔ0v&���z�	�+��&Z�|l�$n7Xu JI�#z5�D�s#x� $�wEh�1�f4�)�o������ɟJCg^�|�5՟g�r��ZMw�3c9`wP�B�F� ��w��krI��r�Z)H���Mx0L�m�T��v�][u�_XKv�)������m���@��:����W�,2m��YD��~
v��,3��g����7A\�^ğ
?G���i:�fOf��ξ+ �x�,����y݅u�$�H�v�||�P�y��z�)�W�b��=?O�?�byX��F�u��}Q�*����آ���T4O�O�9�8�[�{�3�e"�r§���T��}��0U8���z��n����>��P�x�}�c��x$�H�ӔQ��`5b����ޭ#zv�;U��j��j����م�M1e�w!�JW��q���좤8��\y!�����e%�^7�����3fBY��t��1��t�����h0x-��3R�����k���(l�9i$𹈩�T� vb���<Z�f�5fg��H�Y��I�af��~��k���9��}��f.�}�l�(1<;�Ѕ�}�~¨xM�i��TS3���[˨�����!VcGבz 즞C!\.���]����t'4C�%��+�=(1��<	E=���B��w����:M�P/����ΞVi��>�i�����b�TH���G���p���Js���CZ�2�՚k�+���Au�)�±�Κ���}z�<�����qEl��� -_��S��-��.�1�u��4�S2�%�.7?u���&�5f3�շC�7nDt2��2��T��@*r|Yd�z��l
<�]B�L��؄�����������f�3�8�D��yn3$�a�����!r��?���L$�&sޞk��r����7
�������/:��"�Z\!G�}�P5N0�� ��v;@1��u���t�'���� �ذ�Hⵤ���3 �j8�y���Sާ��}R���/sk�$�_;�����ۿ��"͌h��|~7Ig��1�I�	�
.ޖaQq���L؜�}M �։A���>���E