XlxV64EB    7a0c    1a20�������)|��c5y%Pru��S��K @���:1�Kس*TB�k7���w������呼���Y7��6@V����7{>{t�4�h�6�_oF,�<}9"�?c�������t��%5j�Z�q�l�͡��K�i��s����y6+�K��xd^�����Z����=7�o�(`B@���a��}!bH/}�'߱�izD��������ɨC��},y��6�ߩ������#QB��Sm�.�.Я��~�����&cU2~��S�?�mB�J�%�1��W[�K�@k�+;�	�6�#�pt���zf�[\J?�c���#:���;>r�Jį;����v���Q\�����%ȇ{�#:��.�``�����@ᘃ����.�c:���.�ϧ�/fJ������V�:ꚭ��|�<+�rK����N�vN,��⌊�u	�E�sB�0+� hB��u�J:h~�pA�{�J��t��������G,���}7��Y-��+A����P{	`������n�)�y�?�0T� ��W��[��<bQ��w5�[�l2!6����j,5�Ǯ��Փp냰 M�;�\M��%(hq��s��Z����F�j�������B�X�lއ$54�^ʳ{� ���s��e,Ղ��9�o4�;3����
7�� H�~����(2���E9���N���K�˸�Ũ;�R�I�>|.���%�S�1�x��#��*��KC�ȃfm�f4�AW�[���9Np�
�c4���X�*��56�i�@�.O�$ �*�M�����}DUrb9[���on��Zs��م��Q��6���x|�/�k�*���B�У��[�	E��e�3���@�o�H�3�
�:���D����jQ����-���r�$�$� �/G�5�;�"Z����0h97��b�*&��~8sT>B_t9��&�J������&pw��6�8�p^�v�|���||)����p�]���/�D�-v2N^8��;�͎����C�>���(�U2p��a���S��4]�Joic֟w>pCt�1�-9GHe�Z^q������ȱ!e=�/M;�Ax�~T�M�I��y��]�;���g&��%�f�PH%ж�KS=kJ����G&7���q���[<F�����,��1W��k�v��31�
�Q�4����ؼ�� A�љ/��D�Dk`�T�Ȭ��/���8�|�����ؑqOX�g�r�^��cBZ�;�b}��l����̹��U�	m>��u���(�n5��]
���Ή�"�։��{�df/��h���Ҩ�j��ٛ�M���o#�����ڊ���V�b)c��=���--b�Ʃ�e��DSh���4 [��_�O�Zq�u���Sgp�;�b�?��_�~+�r�9V���o���Xi�������f	�/��y�
:�=(�O�Lv�J�zW�
[k��E�Yr��z����:#`�:7�����Ȥ[�x�B~Xl~b6�Х*��F�pCl�'�XO ����_�����ۑ+�̸-�EyGph�h��+Nv���Y�gm/���V?,��C���l��Mӳ}�w2�G���5bҌ�Š�����R����#+.�م�wJg��k��Gm0-�UH[�2���Sj)p#( ��0�58��!>��1y<jN�i2��o����b%���	�7v��hܟd�(����y��B�m9�s�N�L�S�Lٵ�>����`�.B���5P_U��V��)�}�?4��7�`t{�"�C*�dЯd*�N�'����HPc����#-/K���y��3�E��?A�����ڨ�kf�s��ⴗ��-��X��*��G��º
��n|L��C��EM�� �2��K�ײп*bu�Q�A�/��gD�^���?l�Ǿ"���Iʋm������ڒFt,�$���+��g�V�l�	�ƙ�
>HY��wl���@?)��_���1q��{����w)Ye=
��m���壄��Mn��?'�M'���K�L9��[37U�O#Q�*{�d�.U�4h�llC�6^3*�
�Jͅ�uddfm̛&t�	�>�wy������:�7�`���~�_�Ӈw�Xt��ή"S��Fv��C�\�#��N���U���5�9fpEaH�uZq!c,!�.�CK�:�4��1k���@N�C�7�X�zVdv.<��S4�1nF�L'���6��:ʖ�,
&��U�Y|���Τ"(�̇����j��3��cnab�z�������
�2��)�q`�X�)� �b��2q��Eh򞨭(/#��:6��]�x�����QS+���8cj�7�� ��Ef^��Y���+A@��x��n�z���	P�D�}n��p�hq�7�~��<u���i��~AB�cu�u��HT�Ҹ:�v�~�"��b��gV�;tX� 05�S��w��]o�ё�mXPA�x�V�N��u�t��"�k�svrI?T�-�V�r��+;�B(�̖;�ڰAw'��{�H�L�τ�eI�D�Z����x�?I��������M$�;eV\C�)�� �#�Պ��J5A��f�f�l����Fxv�Nc��ئ�O.J�d�L���LƄ�Z81H�}�׍>$̝~G�ef@b�Y�$�62�G4�2��3�r�x�K��R�����P��z�Ǆ�Tv�e�(���5�ҁMb�������I�D$���UC:����K):5n�`��cN�]�
V�dhpB���H�GN�H�$��]j��aV�4z�w� ��?N�@�.3�S�6��k����β�Ή�ܧx9Ъ(��/|��L�2�S�����Z	�}�y��hz5�&�2��_ 1�t$^�'�I���1����A�1Z�:3C��^��m-y�J�]�a*@�^D�0M� w��23��D�v��yu���,ۜk���Q+��Q�$�mP�Aǐ��vA�4?‷Ċ�<�����y��`��&79������},*�R��<�8�n�n�끖�"�%�)f�T؀Y?���̿+y�[�}�.� �2����Gdj��}/�8�O�)�O3#�� �����$�-��X����w�
:=�$Gҟ���"Pg�o͑0F�����(K�6 ȥ�[!�>�`�k�̮�|�j�U�HGm��uB�t�޴�#�Y;e|�W�'E�Mm���']���C�u���R	�ϸ��ͧ�PFI��� S��Z����&D ]2E�E�	��a��0�g�Q�~I�pE������J��L�<��l$��u$_��eAٴ��Cl��i�J4�>p�s���\2��$�� -��`п�꾿!�A*n�3�K��ϖ-Wg! 46��z�i�q\�:�V�P�W=�ϋE�'z��k�W���؀#�P=���I�ő����*�����%��R�	_F�����B�<�;�p%?��c�o�&�@W���uN��<��Rj����O���C�/單�4I'A割1RBa�a�]��_С���Ǽ���u4�0�"f%%I����Jzi<
Յs.�|s���<ķV�*9� -���N��¹�<�1B���'�b���R�>sW(�:64���۩n����a���5Z�t���"��`�b��2:%�[�8"(���1���.�����3f{����c=��=݌��f�|F��������=�TD?�Q��t��jk��h M'ơ¼c�����Ru���
���,a^�.ӓo%�sYv�(���p=%QO��8�Ͳ�*]|ù�������-Ԅ�,#%�����j�-Ҙ+���J�CO�}��E�j��{��1�q���LW�0��tJ�*��k���Yw��嵋���I�R��v.].v�j��S�U2��zyE�s/��D�
�/�i{�$5��8�nS�͈�2�������Ħ�?������ �-��\�r�_z]�s��ۢB#%�-��DL�m���T:}��@��+�Q��%Ns���L�����X�1��,��f����/���|��"�9va�70@Ҝ� ���Z��3�D��̡��̅O�'Q�P��Do�����0?���+Hҟ���6�`ۨ�r$D�T3��4x�I��#FU��1ߩ�Q�H[�I3}`�ٖT�^�7�p閛o>�������w���z����Cr�r ���h�0�g�U�X����x�ls3y�~�]M6N8��ʀc�):�+�QB�TdA�V�`x��Zfq�M�TP�+����X:QH��hV��fW/M�6"qf:W�|0oI��oi�=�����E�)�=��6+vʸ�=�9�L$�#���K�gQ}�Aݮ�sue��;7���:�P��@f�s��.U�E��8�S�j��n�qU����j�w�u�>E'��|3[| 
p�Nxn5�A��-��9͏��8s0a�>����@֡�Q������j7��~�m��Ȟ
T�p^{=N����T5�RnÚ�T�-m�O�#F�*6M>:)@ed�ׯ��,��Ԙ����߽��sY�v���<��V�����&����*��7��>>�vR�$n�<�m��B�,�,|\���+vf�I��Z�A���p쿷Ϗ���D��s�}��a~���/c�rg�hPW�7�������8pȟ!�0�-�,���? '����ML���)E��99!`+�8�;�j�CI�xd��f|����9'G��$����u����a�s�x$��A�`�kV�5)�@N�*Y*�C��-��_W}}#�6f����y���$�N ���m����x,�DC%g�45��I�?���pm�����:ݣia|��8�����"��/k;�	�rw�/U�CɮR��G;r>��x���"��P���2px'�3�G�\�-2���?&f��zD^֋��\?@�s#�,MOy�Հ�¢���b����э�h~I���s�cꧼ���F��?�����K]�T�����O+х���}He�����L&�3C�M����N�s���Rz��+� CD���z��A;t'C�5�)!?��F��$�s
?��K�� M��zg�T8��{W����4�čǰ��_�F�}�M �K�m��L|#o�n��ˣ1�5W�n���4��jixau���>��%}�s�ɒY�*�C�n|���::�ңi�������Uc��%D^>�����'l�ntz��*3���)��w.DN���1���m�0�*#���s�z<�O�eEo��W�;��9Qp�SK9��UE2(h��y_h���N��'-|J��&5L��R����ި��*'b�\��sksQ���%ܮ���M��b���)�R�!Y��i�5�W�^z��]���~���~P���ɨL�u�K����5��b�tC�㏾��`��80~��3������I���^�_8/̶��b��驘�ȏ�p� P�4��e�8h���-���Rh�O�rB>��_��om�¼ @e��,f���?)
T��x�]�T�h�9DI�5�l���1Vǳ�L��Ψ��yp7~k�>�<�?)�� sIx��oa�K����̭�"τ		��j]�[��!I7\�N��Z����1g�r!�/����=�a8��XV_X�/+���-�ǐ�z^9�r����fsc���>�!��ے�%)칪��Bҽ��Ή��Beߊ��ޓ������s�sǼ��)5�-��z�gL��"(�q7���ڇ�m��53Ve���F�ۈA�Z�7�PM�?�ŀ�V�Q"��p���z����FbX�*|-���2A��GoZ��Gy��C��,F�ĕ�&��Oh�_&@i �L��9Pʞ.��Yp��ͬ��D>������m1$I�_�p�?�#���;ڔ�e��Ԯp����������F�%1�^L��ڧ���*�5O/��蓮��C]=�Wk��XI��2�vx9J��C$`�ޱǮ��J6p1���Պt�È��"��+
j��/�H q$��5����ࠢ��yN�ּ����������mU�7[��.BS�I�s���ř�wy�f����~ ��RQ��o�_;��k��s������(5�� �	�E�Sc�j&���������RTz�`(D���	|���A��NZ�f6�֪�պ�=7�
V7N�/����/�L��N�lC��N���<hI�/��4Ʀ��l��(�PV�%=�X�c��P�Ga�a����0@���Ey
��|�RCJ�X�����f���a�[ZJ#��;�3�q�li�L^��]��K,����MX�xc�p�o_N��lvL�V@VN�P�k���;��\��Q�5^�|B?�V��n������ۓn��������h*=����ѱh��ρ~7�����@��i�B\��4�3��:�7Y�$f�{��XH�Qϻ�nA8Y����`���7O�Qצ��9޽��uȇ���Hf����B3߳VH ���	����`Jq(��t��+��J�Nf�(?�����՜��@A�W�+�����BG����M�n1��M��:v�F�@��lT $Y��A���W�355G��c�o�td��&��q�'���k��@���H�5`��L�K;�,��<�" �w:�W�M�N�!�m�WA#y��>P#������\=�ÐL�nm3�