XlxV64EB    726a    1750�l,����om�]��<��xb0�yxm!_eC��h*���ѫ�~Y��?�U�Ƹ�ㅦ88�?�&x�,���w-���57�� �g�M��;�	��V׼�K�Y �R�'�rL���
���n��Y������,���*�I�fy8d�b��DGF��I3����/S�t%�ԫU! aH)z{�kՎjD�QR��KK�P�Z�Z����U����TO�m�������n�cfe�!�� �j��cd>�F� Q8��p���!���$���?�pq�{���nsD�02F�pd�k�Yv���|$m}�Q5�ѢJ������D/٤�&� ̀�/'hV���F��.K��vo
�WZ�q���-��/��گ��~Y��c�#��=RGO{��wّ�}^�
�U���;?ޤo{��g�z��i3��0�������j���Z�`���\���s��K4<��o]_
�n͕G��PO��Xb`����2��5�-G�N�|lX���l~�Qc^��Ei�x ��ۧN�鷾X`A�H�ш���Mŗ�ͧ��x���E���@]46�_qx)�ɰMO�.�_y����mB�Dc5
�GP=��.�{`�od�xGC���P����KOp`UgdD��ȑ>�2��ŅK���o�7��@L6qO�����Ti�cdW@�ـ���ew�`>s�ЙGb^qH�}6��G'�-a�ύu���m:,܂+I?�j��@W�׽�O�~��U���o���t��î$j�; ��m㲤J3ΰ�VL����^��ҌDsBҿ�iq{"�JlC�Sw(��69�e#���)��BQh0�a�⋭���/����iUXL*j�5��	�=.�i�tщ7��:�X@/C�ߨ�Gƒ�p����Ό^h��y�� �K��dg��b9���PʲƩƷ�~w�=�<_��.�U����߃�,����=�l��o�c����.�0T3t�~i�JŰ������`�@�6���{�޺��?Y�~�l�DC���F�UUa1VP����Qd���8y��y��jz�q���\�r��o�4�����!�H�r�"H~���2�o"��;����	B�@B���}2}x�P�����F JP��"��}�r�/"���>W9q�\9��R7N9��y��hv��0�:����G�- g�����:RT��ڠ���,�]�6��ǎ��y���,~<j6��������)�a�^��ʁ��e{��M�J�}ܐ��)3�yb�\��]�sb��P��UN3n�t��3����r��M�v���C���&�s��������N8E2m"���:��� ��72��.��/�on����@��"���ܦ�;yW݆~�?���q!D���H�nz�I~5cr���2�^���Ǵ���㳄��CY�<&��:Z��+G&>@|sMLV����f�<Oiԃ̫�
Z��6"�������Y���������:�d��N4����c>��CV�se��98���U;�����-'%c�������6憅�j�?(�IZ���1���q#�K�Jc�+�oM�J����w�x�A�n���aA�T��Ć02O5g�}�.�>���������o�c�*�K�/�G��7K'��V&�w�:�0��;����9a�T.�o�P;�;(J��IXh�
�Ƌ'��w*��&c��_��4,)���9��3V0�1��O��{�B'�+5��p_�w0e'o+�4���E@�0\::;�ȇ7x��4b�p�2�s������H��^�}���Fj�USO�k�9ŜE�/��<h?z@�8�e�#$���(B�C=Ն����R�����`��ಞ��BY|��,�	v���Dy�ѩL�!�4	HU�<�\Y����B�{<��LXP���s������n����0�V?���;����X�f؇��1�����4?\�����y��p%'�뗯'i���M�,M+�D���sQ���'s�_��0&�1ҫ����^w�>�3�����NNʄ��*Oy��rO�<r�>��K<L�!�JѦ�쯲W�g�*�GK�k��L2�%�2�yj�?*�`sNcT0�(3>i�>�ԭ�.4c�i�o^'�=J�M�`����'&�ܴ2�_Ø�x*}�9�dN�,^�hSQ�f_C��񎷎C˴��_Z��CNT�Ch:���&nF;�8�˽1���B�Jqi�.yp��^KO	r��$��	���4��v�5I%>X����lt�3�~��y�WH�����]}�릏6�Dtu{\�������+�E���!#JA���Y	�sW�ӧ�Q,��t���L�.���#���0+�%��{e;Lj�rQ�pݱ��4��R�7Li�G�PJe*�do�e�z���&Q�F��Q�/s������7�f3��ͥ:������ڄ��Fi]�@����%�_Y�Y���w
0�t �]��	RTXC���fi�-4} �LT�sU�EwO��T��bܮw��� ��SL6�J6
��;�nN�x�N��&e&�Uu���7&�{SGwsn#�F&�2�M�u���� [Oй�Z$}4�g�f���y�����
2�@$�3ޚ�3���sxL�#��7��>0Ǭ&�2�����t�Eo�eƎ�XϼV�� 7:�^�M�������$4�f�����P
h�,p������'�C8v�˨-#%߬� zh��]�F���HU8��u����ܢ�v�c�@˲��4�rP�]n]��B�{�xǅ�� V5,��\|��|�?,��u|�����L�$RcC<���{��R{�9Ev��VF����g����"\�S�J �懲zu=���C{3Ww�����@:�ɏB�N���2@d	O&i/U_�]��G �s
�$�Z��G�!�5����/�t-ħ��a�ԏ��Mz$!��X�h����Σ<O��������#iB�8z'u3. ��%g�Ec� ��HXvT�T:��i@�t�#�!%���~���§��\��!`v�]��T)f	~�ݵ����ހ���K��<�����i[����+Ncv,�]
��@"���5�p;'���q6�N�n�QRċ'U9Y�j�D�4�W���tz�g�)��Xn9-���P7�ڠC�&�˺�
g�U^��U�'Z3�z��v�낕�ojvT�x8��ci(TaI�C�
�!�FK���'\:[i3W$er�3�5�30�b�#-8RNP�]Y*Ƕ�&�]���~�@��	��	+w��x�$l�e���>?�����Q7aN��=�>-�e��VR�ܴ��<
���ܪ��C���{�6�;��ի@���b=By;`�qӵ����.q̈́�Q�uv�L����|���X�/�+��Ѝ�:�nQ�����-kv�
�K�a|ub�w���'�Λ�sǪ�Q����q���U�I�WE�l�UOv����Dė6�')8,��}�=��zIpaq�TC�ħ�($�z���K��8��I�[��.<��JtD�ӐG�%�rhNL�QiqN�4H1����V����.��G�81q��Lr��jL�� ��z��f�5��E�5
@O�<2�b�4�.%W��}�^<WW �Q�[�S�����(Bn�S�)2m"[�To��o���֐Xa���h�k�Ŏ�"��E7�,���)�_��Oڮ>��B�p"?:�^���!�Οpq7T9f��q1�\IO��*z B�esH֪#���q�u� ׁ�ڗ�U�+�� �P�V����Y�h�P�XN�PWb�I�18�����B�9���`z�3����X�wl3m�QO���͒��r̥��� ��ꆓ��G�J��&�c��
j�g.��E.=��:cDH�b%��b}6�*X�w_|g/A�)M��m��QQ��������7:����E�@������3^�/����~ҹ�� ���߈q����Pؔ|�^�1��68���m.qc)3��6���=�ڶ�8+C�������8�-�fpnV�F'dAR���w^^ L��I+Q�k<�q1�>*��Q��[K�S�mf�����ʃ�}�(�n��� �Էq-�7@c������+�ϴ�L�~��YY�2QAV�uT�i�J)i�2�w�S��i��$CQ����T�#|��v' Fbp��n��"��ޜ+ݳ)L�����I1i0�S@�B�r<�����R�E%�u�F�jذ ��\��m۫V@Ly��
��������g�}_3�f��d^i�K��M���|�l���C�z��f�*��.�{`
#ȏ0����[#�@��i]� >�FY�޷�`%t�D���	����C�
��A�[Lv�[,��~�3K��L�#�2����@��s:�I�G�H�t��-��fl����"3)�a;��Ԇ� �DĹ����Y{1&ߡ.+.Jz�9��؛�6���*��{B��
���2�"<XWq�wy.!OI�F�g1�#�Dr@P��ѭ��c��p������!�k�n�\�2ؙu���ı�֬�s%I4�Ipj� ��B���U܇�,I��]
G��gr<V�k�!(�l�;HV�7��p�'�`u��&8�����4
Xl���Μ��P��.�;0k;[Y�J=`�`� &f_v�diFn6�Mڰ�w�nI�H��ܩZ�8,��BF�����XA�M��9����8_i�l^|��}1����M��/�ٿ��:��R�A5�v �yj�𻟆纮�6��^=�$Xz4����7,s=�<��bf�n"Dn�]��'S��V�8�������� Uic�_N�k��KLٵU�2��Uw~�0��$���X�v�� ��*Y'��v�c��܁o�!W��9��T�3���yT�lG	Z����8ufӮd&P>���^?���yC��	��,��lP�ɍ��\x0찪ty��q��х�fpw�1	gf�됥�:��aI&�}�C��-b?�_��hM�	�!z�*Z�vɄ���� �<� ��t���ԇ���!�V���|��y.�x������ ;���+��D���Q��ڔ5��ZIL�zH�#$�ej�-TaD1!L���z��u���Wq��q��?�R@�Ę�n*�)�_��U6^��/�0��	��X�P������߃��	����+�#G\��v��B���|��H.�@�� G�`|{b����	��ho�#�/`���__��je�����QR:�ฉ���NÌ���`c�lf9����5�q���2A������4�ڃ�:�kfy��k����\h��yo�7z'oU�rg0��	?t����+�7'q�a�xƗ�I��bMo~ ��u�po}Tf��'������}� g������M��^���Y�m����!V]�v�^�:MT (n/�\P��������e��{W�v�GSS9Y.`gGx�d6[��8N���i��;��y��x�!��#��T%�JTt��as������֭!)n�.�4�M&R#Y�b��(���<�������c7K2��� �R3ў(l�(���1K���BkU򖱶�gh����F�4b��2�oT߲̘̚9N�d�J�e�s�cO�����47�s��c�4��k�����O�����T�6V�9ӽ�ΪoS�0�̽�v�D;}���,��F�r�5�4l�����g-�͢M��w��z�g7%��~��6��E	^���T��`����>�C���J]�މ߃-�vMS�z�� '�ry�_ad�3�[x�CMk�Õr$#l���gL����
�ʟ�,�dZ[�y]�|7��(|/"������J��D��eyf~�{�~�sx�0=z@M���p
f�SX��L>���6T�mZ���Du����D h��
`��s\i�E+�