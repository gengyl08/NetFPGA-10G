XlxV64EB    517b    1220@����<�qX�;z��h����;��>�s
��7�����O��?���Q[�������YP5�����m;�aH�0"�v�9;�`�63HU�f
]1b�HH3j�D�ބ�]Es-k(0�Z����M0���zG(�Yl�f$L�ص�_:���f�9z�UC��I0�%�=h����~�".�M1h�}!�i�To!lɥ�Oq�E��l�U_RC	N�?�e95��
#��I�2"�T`w.�=��(�#�+����l8MFD��d�����"7�5ҏ3�PymY4��a��|fB�O�/���al%	��M�NO[M����"�J`�MX�Q8:��蹥��b��� I4���Gw�����$�(_!sl#^�)��|�O��;/�IIe���ͽfm�#˸}'3'�F,rף�o�Ʉ�|B������{�z������})�-c^;�Ľ��h*���_�#�����(��B/��J��E��HZ��
u�POP�/2��R�3�pxc�"��P@i
i-H��&���گ�%�l�l�
�킬*�X
��L�wżXB3@)O/���'����¬���p����N� U!�&��V�E���XO�c~+y�.��8���T-i�S6��Zx�����	���`�b���B:O@��`2�*^�<�����V�yQ>��$��/�"��9�c%;���R�}#���W��:�P
-6y��jw�H�?j�c�'��W��P��@k���S�Q�q[Z8�o.R&BI��'C����p������Q\�G�_f�]���Ѕ��N���}�]��r0
;	O��K�����\�`�j���Z�J��`�TM��Poz�ಭ�G�d������Ԁ�(M}Ŵ��� ���������w��P�>E,4�Y�[fm۽���$�T�|������j�,,�փ帄�o_p����?7m���5~�;d��_�|J�I�
�f �ZYfj�Xv��f�(	2�˫-��1�*��&����Eڸ��hjN���W��Q��t雪�����w��@`n�����;���*tS�X4��I(��@�;p�x?^��U-G���Cd�듏\�~������7j�r�h������I�[+��	mA����06����S�"MJ�Ã�1��	N�$h.���.��Jh�g���4 @,HU;��d��p�A�g���S���-�ـM#ü#��߿��=]��0���odH�k��q�fHhg�u�k|O
5��r(���rG/��Dz7��3��}o2,'#u"�<ns��H_:��$v��K���&M3�%�Ro�64,��>�zW�]�=X�̡%X_��hډ�W�5 h����FWn�s��5�B��|K��a�?��~y�P@�)�
��x��5X���?0�ZC;u����,�S?־��%�J�ѥ�ԓ���@�W��������8^����J������	�����w�^{��O#�J�q����ڏ�%1�!��F����n��!��l�ݾY"����J�n�*SJ̫m�>�)�D�0�n�vQ>���7���&$ˢY+'��6$��y�t�vzoE7�(M&^�������T�\)Ri�<�S/
�F<�m^�&�Go��~0MMhl�D��2c�=U-�d�f��}3�M�9">.��3 ۠~�T��������{y�Ow� Vf�=���aG��_��HV��)���� �������-� ���K�'N����1�<R�vG�i3�ρ���}{�>E�kq{d�|o��#ł���.����T��@�Z��{2H��B=�wQs�j�x���Cd�z�2A��g�z3t��i�ѭ�wk��ZlH���w���O3ٞeI�`�7H��C����
�k�~�Z��#May�6����N1	��l�ҩbyiNϪ��ټx_�G�� )�}ȏ'��Z��LO
���Pm>ݧ��V�Qwj(%�[A9���1�.�;�1�@w�,s��o�Д�	�>E��C��w��޻`���}ZN�E4��z�&�6��1hk2I2�m3=���9b�I�0����\�з�Å���{�q�r��Z��N:G>4�P��j%N(&j �C̟g��>���AC��8��7�`���лlؠ:���aj^��=���Ĳ�oL^�-����z:p&�"���~�?�T9����^b�Xr���|�`�y6e-������Z��9҇#�r�n8Gk�@!��jM-<���\4$��'��g`��P�Q�`��%(��P��K	������{%�η�7�Sua��U[�)x���8ń0�L�Z�`	���1!���CYf?oc��@����Ä|\<7(�:��/��c�Ġ�� ZA9�~3�"�ȯ���jN!�C,�,�U�2%de�f��M�X]�&`�.H(�p�$u���u/�!����f��%�;v�p|$)rڲ;��A�WM�6������a	���E�l�|�w�~��~ ���j�[l��`�M_`4�,+#��i�q_?s�N�{aW"��af�%�P���wo�yk5U3H�˿�r��j�7�5���5;R�;��=�Ű3=^��Y�Q�$�6�>4�	����~�jaǾh�z^�u�tI�_^����D���T�*��[y�h��sx��u�RF�X�˛�L���ˢt춰�Q�Ro�vX���^>cH4eG��ź�ô��~VLv�������0�'e�>�h㒕�Z�`���Ƒ&��	?�HB��V�4.E�q�J��?�szI363�5)�� >d��q��{e��F�ɱ��R��.jV�u��Q`�:2e�v�e��u����ICJ�:M4j��A�9o<J?�K}�r��or SѺK���i��7��y�	t�JYG���M��"�N�8NM��܇�iK��q�~���	�=������,�|H;�Jy9��7Ě>��<.C���pZ��i�� ��i�V����I��x��� ��N���*ר7�rHfZ�@�IKy�c{=�b�y��x�����N���.�+�q4rt�a3���Yf3���y�S#�K���c�H�u��n�{��[ݩ4�e�E���4��g�&�2����ia*��`5[I���W�wy� L�û(�}�07?��½~��_ԣL�gioAY:�T^Uǝ�$�[nK�`��z�|��8�~u�!�~�n�EI�ŋ>�W:�,¸<��u����,(3߮3��R�8�RqA����+��a�Gʼ�
�R(J$?S���*��%���K�B���B$����$�+պ�X��"	�饧T��G�v0_r����z���K��=�ĵunG{�w��Sw�iR#�����3��Z�t�	R�x��-��w��L���z<���v �(��Ծ͹��H�vb�vF������K̚8���	�n�=b��&M����@���_��ww���BWw�e�d�S�Ӂ>-b�|��꽣�%��j�%��(�"�����;��;=�������A���;x���f����܂������}���]��Ա���Ӧ����iD]]!mn��ẕ�ʭK�^��5��aE�Z��>��|�+�D\h&��o�7�������0�]��7�}��.mm��:����W��^��w4VU�����5��*K����G#ӹ7u�ܭB,!֜ȹ0������d�&��`):�����-�KH�m:�&�����*���9�r���q��c�|"D/"�'�˛@k��i���@�F�B]�C�_�Oz�s<w} VNV;�tP�#a�n��rs����W���Q������V���,��2��n �)
V�l:�G:��p�	?����(�Ԛ��P��v1	�q�@i�^<�&���v�46u��r�;woB�^�I1+t��o˽�kǪ��|�WpO��������h��O��Ƚ�s�~kk�ev��Z���T��Z�Eq$Q�p$%���흵\~��7[�,���S�����[���.�QH5F�-02���XƏx9�x�)��R��?��!������j�q���i̍��]���{v�6�'�`@3���d[1�[߭o�qD���R| s+����,��3�\;� ��2���r!{
'�4Bv��k��Î�â}Q�A�� b��a�p����uF/�a��q�4=�ʆ$!U0v�s:Oq1�����p��HM>@T��K��J�GbC#  -9W:��%�H�|_@#���q���j@�b��{�.ƌz�9�ӑȶQ"�߸�� [�[ ��DN����T�}��a��k�wqƓos�*̷�g��fK?oH$<p�Ӈ����b�.�2d>�yо�=%X���%��X��E��֐3�=���wQ��T�CS��B�a��j�"�C^��ۉC�=z�,��VT�2�B�v_�@��|�Ru��j#H��#9Q��H1�_'�}�i���+�w�j\ �:EX�~���."TM�o�8LX���̩7K�g�%�]OO�LōEg5?1�uw��x��F��p&�V��S|V(Y���K��U�ro���jÅ;�N-���r%e��|Z�q���Pt������e�q�8�Z ���@�X��1