XlxV64EB    249d     c60a��p\���3!���
�>{�0��a�+C��|*>׶�۲X�ڐ^>W�vO�#��G:�3��B&��v����F'ln�����ǳ�OP�{
���^�4ҿ(2�5:bZ�i�ݼ�5�y��5M�|�'�wl�����*zjxbz
ox��@+��a��'v2r��r�t]ĥ�x���[נM±ǰpV4��!W#�}�KG�i�`o�{� �:�Q��x�|���r�`�	 �)�-��j�^��1�Ŭ�|��!�E�[�r��B���_1�ZBB���	�b��U&1 3������PMn�YƘ��F�*�F�K�"����QRQ �@oo1;i��o���#h��r"����e�C박��Nbg�=J~^�!(.��(��k-9��0)f?�����|����]�z��Q.U@�*�Պ�0 B��@Q�B�Y�aⓓц��W��t��X�.1�6o��v`10[���?��X� ��}co��$O��^J�O�斋���Ѐ=��ЭΚR�:	���͂���W\*ߴ�ԃE=:g���.�-�b���<����饗_j�T�LGޯ�/��4>�C.}ьs'�h��bn�w�#/9��eS����/�����W?�	�_�־���nDlC��!L�T��w��_�%|�(�tڀC���4<��ŷ��5C�fML�W�kt~�Y�'���Y v9�"R�y�����Kf':(���Z�.�Wb��!^�ʌPd�v����U\�%�`�d͘c5�)P״'��8�Z��+�?���t��3V ;��KH}t�j����ߗ [��5�0Pr'@�H�ˣ֟苫��襙L�x�XP���,G Rd보:��h��J����n�C��E|��{�+�wM��'�o��4.(�5+hZ���B�6�Y��]��PB��y�Q�X�����_V�k}�Ck�+��tP�]��&��zø�˴mǝ�`��/z���7:ӧo�ezx���������w����'���s����V�x���N�����8#y{m���E ���8Ǯ���>�fA?�B�ʶ嗐�"���@�G�~�%vJ��4���,"j[��.�i��� ����wՕ�4|�O%�M}
s��q�ra�bd�
�wjo�ƕ<ֿ�C�F�nX:C1|����Էi�)Q��'h?�Їv*�ķ�z��	i)g9v��ۃ$�ӳ�omu4�؂s�Z�c�6�$�=��tٲ�W[e!0�� �y�n&݆>�v�U�����N����R c�f�.;yp�̥b��-��/�2N���V���~��քk{��w˂�T�t��JzrL�o��빦D?H�~>r�-r�;��
�*�r����}�Jڹ����Ԯt����-���ɦ����|�1��^R�oEm�r֘�`��)e�> �o���#;�/* �R&y�>8��*r`�|���^�����֞!,X��{���ENOdՔ��ڶ�`�QX>s��J�L�6` "�K���<���T�ތ��LFн���4펣S�FJ`-��t����WBx�jCو��Q��_
෱��*H�)��|'Z��;��m�FɃ��J�|�?\�ճ6n6$
��������@�}�'��L"�&�p�Fɝ�]}�!}1�T�:��v�_���v����:���d-Dѡ�ܷM�Ҡ]M���;�>k�	���\*|BG_�Ȑ>4Cd�ڰ�	 P�Jl���]��M7̕�Q�~5�V43�!Tn�6�&��-G�1I]�is�����B�ֳ�G�vet�%���(�UZ8�I"=����!P�	������K�R?⯌��(`E%7��2�46j{[��$��TSx"�?C:O����:����\�kM&e�~ �u��nM��7 =*'�0��!�zqa�~��K�5��-@�JV�].gb��4���|)؟y�@|���u���;� V�&�$��ܜG�	�0�A�ȸ�[<�)�b��2��rX����������Q �:6��)�{%���=2査[e�n���
�XϳU=U�Bq��v^A]G"�m0��|��ֳuȵ>/J�i�8�̆��V4�ݲ�e���q�F8w�2�F��<=+A9~����լv	�&�s��m���F3<<�^��;�]תqu�q��2�#n�� ��∆,�F���|�׆�3��œ����>׿�E�Ǩo�O 9�פ��!�VaUMR�PB�Z��ֽ���7&n4����r(��P]h\W������!D{�0	7��jC;b+�l�c�YC��=C��<E�d�����Ԝ��[��4M\��`ͩ�-
�1p+��a�t���W�Hx������ �e ���[A�@]�?���H]�d�Ҋ=sA(�c����ZF��k��L�]0g�S$:h+@����6>]��UY{y-�U����qX$#�2T�M�%��w(d��+F�����9Lg�Zf7af&��R����6�(zGo���}�[�=1�(����]��K�?�K���`���`B�)�|�����ՓpO� �C��E��@�P�\ޣ_' �B�&%�aA��^��L���x��'n(��z/?��L��:�ͻ����pQ����M�Ԟ�І[�������fm�5��T�мL��������p�&�#��W�ݤƅ����@��Z���w��^�� ����n$c�h��j_K���	�����Ne���
:4�,=��U4O��a����%矞[��E�T������s��]�d��뉂q_����~̸a�w��ukG��(�u{�=��k��IS����"�'���O �W�(��K��+dNO9c��o)���:l�^	f4����{�a, �����W�/0�
�&feH���?eM��T�v.�� �W��O�=��={��5�(�7ϓ@ E�V�$( �ʵV��jI�y9}aoñ1������w�����$���VB�#]Hr��1'4�$��B�;a�b��t�>����������X�Q�);���\��dw���jL`xnU �|��~ҽ�;�Z���\�9�KX��C��h0�я?� ���=�yw��m��J�d�S�v�P�9C?}�C_��;5Lυ[b
���b�8��]/���ƾ����Ǟ��,�