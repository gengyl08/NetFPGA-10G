XlxV64EB    1945     9b0�F;�\""K�����z�Ɲ�b�q�u���tW�5Q�]����wb��K]�{Ǹ ��;�3��e��j=�P5��
��M���P��ߜ��;�쓢�g�=`���g��Q$���E�ř�i�S�*�Ӷ��Ȉ�%�0�D�h�����)e9,�+�t=�dd�x���qq>��F��b��r�c�/���|�Z+���6��2 �����dӬ}��(�4'������|�e���I2���\�Y�彀ӣ��Jς%��k��<]��+0Y�/��@�a_.��W���q7�P��_Q����Q����ŚA�~�e�I�p�3���Yl�5�b������;�.�隀8�~�tIf)�i	�{��dMSG
�"8˃Ua���Ƙ2�/z�ycˉўG�Dv0?@�&�N�9*"�,��i����']�M�[bvr�.Z��J��`���9�%z_�o3{�QPԣ]��

�E��5��0x�qO��W���$R]�Px!΄nٛ�,�CqW���&��Y>�4Z6Ozmບ�n�
|�5��l�'ftn��$��	B��$*`�VB:����sT���p?��Q>�a_~}^��`M<�	��#�]}.h�Ln����&�Y
L',~G��$��K�����eM��u�X'�F�70\o#��[�\#�IeaE��s���%� �q�|d�x���wk�.tz�ﮝ��h0p��gy �4�@��Ͼ���/�b�|.��u��x��14_�:���B2��.�i3<"��K���ߗ�<`YX��T�G��d'#Iփ\��R�o	�B�Z���Vj���0jc7�N�(j���O����:��m!�ӓ��ωD�Cu@#[T���C9(7����\�e���ADKjb�9�Q�3w��*!��dG�=g9�����\`��A��v��V�ː(".z�Roo�%� Q|` !y>�������
�-��r���-�;��2�No���������W zĊ�̀��{�(�ܫ?~����	���O��S���(����$8�tG~@!c���k��*P�DN{�p.��*��mq��'ǩ��5x)r�����-0��Y��w|����7]�ƃy��U�l�V�E���/_9<����4�	J^������O��,��F���zC�R��%1!�W��b���ر�2x{"��<�5��>�H��#n�v�/�����K
�C�{/W?��Lvu��o��d��!Ek3F`�rյ<6��C)VU. D�/	�A���p�� �V n�uYD�х�f"�,y}���� ����%�b����"8p\
�2������� ��k�\�Շ���:~��ky��Ѷ��V>o�f�K����]�U"�Yv��9����p'��`�B4	7�:VvB������mp+Gtx��C�����TS�q����HU�2�{����O3�h�Q-���M�K��_�����&�:.��x��)�ln�_���_j"�Y���$K�>���Z��_�y�����c���}6�0q>
�����hi��S+�S���W��œ�٪o�k�ıl�v
�ꡐ)f4P�`�2�-�Ρ�:����w�����o���x!݌W�aV90:16κ!ri1F#��<�W�Z��c����p2��)���o�c� ��"*bD	����!�)���fHG<D%a`�je!X��8O=�?�!O��B�H'���FY�WB��nMw�ů��2/E����=7���?�$g�Sq��-�F��	��ݺ���5��N_p	����ͦs�SX�6��w��WX�9M��BIz3
:��n�����F�	l�V���(,�lT�����Hq��,Q�>�S8ad�`]�h��h)�7���W�?E�G������x������#}^$=.�1x��	�'��FSߨ�^�7G����/�^K`b˿�+x헪C��պ�u�-�.���I��>Ok��%�'{���F�׎�8��J�vQ_R�5�"v]>����,ӄ&F�\��2`33��l*I����O�Ǭ���<I�ōC���n����x�N_Ы�ZHk��:��.��T9�f�,�R�	�����U��=W0�U��t��~���~ڮ���n�x<�Q�V�c�ҝ�hA���J�M�g�͎�XՁb�)�I-_�b2�>�L�(7+��a�Ŀ�:e!����ϰTf����;��W���,��=�����1�J&�&�[��`�oG���!0߶�����T�����/R�I.���={ɶ7�e?��'I["������XEv���%��9��kC�"�	C���F�C(��u�oa�ʎ>L�\�̕F��Q�W��{�HW�p���3O�/E:�b�:i��������-:��,�q�����V�>c��;h�
�-�*��f�#!ծ+���]��z�����
��?�