XlxV64EB    59c9    1410ve
�E�����}���B���H�;Äo���d���d]ԁ�]�,@�R���ɒ�K��[󑓝پhL��G�>���"#���8"?v&y��~��kG�?�v��J֒��+��ͮ�@,�#1�z��@Ay	F끉��iړ�B�/��cPJ�����饗����|Wh�v(|�3!���
Ԁ�?dO�	�.&rǊ�(�.-ģQ���sX��Y�Ck���-8،}ұڎ5���q7��^J�7Q2CPA:�����.�k���)��"�4G�
x��A�a;��-�]�����&5~�����c=�K�%�S����^� �wk��'B��0��4h�:�a�cpN�N�6�N!�h�'��;�>�Lfi��b���K	;vD��h(�G����s,�ٳ�2�+�Fr�a"��(;�|���^_��h�8�Y�;�Ǫ h���	n���ȋʉ8ZG��7��~vNLR��L9E�d�ƹXR�>�.o/A�؀�"���J�����-��v[�9���B�ƚ%���pIϠ.6X l��p����Q��6t��h�D��� ��T!c|#���eo#[�h�1<&�Uyc2�h�ο�;K@�945�l�
oZ�uq�ݎ-�d(U0���B�6��o§֢8t�7��%��?קO:�r�-���S)����i"ћ�2!x[D��	��V#�jh�9�o��T�PG��9���i-�|{�h��=�����F�[]8j�r4y�aҋ�A�b����Ҍ7������n����-v�Ϭg�� ���Q����y�P�	���;]�3(��0v���!?�>��5��	tNI���P�Q��h
O�q�[35 --펏�j�V�"h:�:�����X}E=�2U橥wإH��!� &�K.�v�/W E�u��Yf��Y " �����4�1 ���x�!�>�r��33��/}�`���l�l��p�p���"�JI�}ؾ�ƹ/���i�2���t�֖��7 �V���`��+F@87f^ݛ�:��b�$r'�I�*���-�n����^���Ǧ��)�&wc�m#Q��5T�.��I�l1$*6�Q�1�EI�.��o1��O��)
�OƉ��5\�YBX�)M�
q����+����q� f�5rJ�4�>�+���"��c���y;"�n�!udT����^l����
ZP�S-=SM Kg��ya�v=��է|����˥&oY����i*�g�HV2j��g��0��~e%ĸ��ˑ���0:�QI�h���c���c��"$�!�p[��U��}]=j�T��(5��2~��NP��5b����&��K�B��X�A}bDޯ�s&���:��jݻ&�����My筒���jڣT��>�_���a�2]Q�%F&��,�%���ւ�f���j���D9zSQ>Ow��Q�ؖ,���L�;�q>^c�U�s���i&N��m�P�R�|f煱o��>V���[�"f/G�C筈'Ӓ
{�Z�Ƿ��-.�8LNb����;��"w����2=b��#:�-ʮW��2��/����a����5,�S�	��D���� ���o�2#�e�!U57#�����bV�oY�V���\�N6�_;��B�G��֊1K`.y-��d� �ř��5���D�A�u�����1�Ƞj�����[4�_�a޾ƈ��<ef���^��#�Hūb��f�/	��`���= �\[#}�X<%�BS��UJ��'(�C��,���<A�p���N��Ƞ��Tq���N�-|��~F��q�ҧ�[��v�"ۯC�#��X�*��0�6ԂL)_[��UE��X����� >��Fm%�[H�B�?��ؠ�X��'/���|�����@R�9[C�O�����[1^�b�3�ƺ��C��!Ce��@�ϫ�j���t�za�7^����^����$ mc��h$�Ʊ�"�� � eZ7I`W�m�o>��I�B���"-(@Gw�"Xh�q�� �q= ���� �
�	K����M��^��DfR���L]����-�`��	�g�P�2�SH�9^-�Ēw��2�O�dib�:T&J^�S)&yC��QƓo�/�5��3F��*�(�1'N�����"Us;��k:���v�@�_���@�$����L�-��Pظ/��v}ᇂ �(��G�L�wZ}Z,�75�!Ac�ɿ	\S�ayy�9AοqS�ν�-g�R����[x����@�T�z���� ]a".��)���H= �qL^�M!����9)�w�#�*\�{�����͝�4�A?�G�T�KP6�żt����j.�����1W�]�rű����������G�� N�,����!�������^R�䶘��rn��+������z�$�l�7"{���g���颗��/�s�U���Ye�x��ݲ��戌V)�
�W��!�$��CL�Ez����B���@�S_l�Tkn�C�_+Z3��9�����ZE+���k�����]�v���Iv��6ɞ;3n�6��Icow��Ìo����`[b��1,.ȵ�Y� o�B�ל�9���qs��+��H]d��i3,���������eY�:�ֿJ(��;Х<����W��?��P�v�\x�G?��Syr�,0��j���f.ti_�n����%y�q�`\�*�M��w�y�;֡ڈȡ\]��s*ξ^H���K��<�z8K��%e���5r���CW9���/V�U��R��Ou��k��@XY5a�'H��y=�T�b5�}w�#�3�$�����=�.�?�/r��_�\$��-��|i�Ulk��G��j��:�7!,s��?��ǟnKlNp��b���	�נ��:�m��
�a�BEs��=ʈ��x���RWN�|DM����\.v����:vm]�"�׌�
0�J���
ٯ@���%
�A������˼pd�l�H��������:a�'����+7b�(qԇ���7��d.2��D/`I^�-��cVf����.gi"y	��� w�ݥ#�]�4@����J����Ԝ���B��p>��1������%�%�Y����X
�̿�\d}Uډ�Y}��Nh{�;����3��1���3�R%f��1t�{%9ϥ疃R��s��w΂-A����]�iXIT�G,r��o^Ra��P|$b���[�I��m	�QA/$��.[�Y��D����8����]`���Rŝ��ߥ���<�II[ds�ʉë���n�$��ܕe�(��7��~�����%������>���%�+qضV��[#W�;2jU}��?MG��e���¢f�\�ϑWm�НI(oA<��'~����Z��r�H��+���y�I��>M��")�`1(F�(�����Lz�b�3�}��vC�dA#`�H�*h�H!Xu��"��#6ib`�2���C�� �W�0����D	���f'�������p��1z����tJ ��e��ZG	>��\����%��t#��ޤT�v�}�VK'1�#�TЃ�		3�xiQ��MW�9�K< u���������e��AƔ����c�����LilK���ʓ7W�yq�x:�%���+^�1�gB���u�M����۸	�~�:"$�*sQx5����Ma�N�en���l4K��{��(s<�����9^4̍� )74-#_�>L� �d!�����zR����40;�T���{&�+���Q�юY`�ų4� }Z�L_9~�p�TV�`T_�(gi��X�@+-F}
��G������X+�IiS��0�Sà�<�)��@��^�:�#�~LUka c*�]��&8	�Yd�t�VG&��#7���8�5��-�����L8i�L�����Xa���0?�n�.�j G� ����Mc^�'�p�)g��n�g�����g�I��0ؔ�n�D�aWK֦�b�O\��؆0�y2IҨ�BSi�_~�m@@��O�g�:�]p(�����z;��>Œ#N�:�h
x����c�����I�>���:�_ah�������틓�4��\.�?RF�dr�l,Na�o�տ�Q�>�%�c6���:���X�US��cI�-����`�T�Q��:��I�z(�l�廛*��y���\�o|�P9`Ŗ��n�����b�2��( �/�{
)Qń� �����ݬ���+O��D)(3��jf٫:��ߟ��x`�'AA�q�/P4'?Gl?]�i�mݪK�T��[o�`�a���x�x
W�3܆��������ꗲ�a�:�g�g5;Q$L����-��0.��{煢鴱5A�
9{��v'T��8I���d�[�G�S�����I�Y�ŋ��*�Is|3g�fЃ�̉�0	j��W3�V��k�.��������B��xfϊ���n�o�z�sY�R357+�%K�v���eKoc�Fd�/�2�_̬.	�[����0���C�����p��5ⓤn�2+A�q������X��a~�׼8c�����;ܸ�b���| d`�W��#?
�&�u��0�t��_u�(����\�K�p!S���j\.طR�꫗	A��G/騒o��]�)�EÅ��vJ�5��Y���	���ᗷj���ӷ�DMf�'#��r#�=y0n{�4��D�>5�ZY]���i3aSc@�������ף?	��5������Ow�,4���U�)-�ʎc�]�=í��螪(r,l?ȓ@������-j4Qq��(2y�SG��.`ǫA)�qG���s��]&�mqo��j��>����ʃmS��*�-�K�ު�NW/�U��X��fB%* q��-�i��U������i�Y��/>8� 	D�	u����N��na������Ty톴���@}����9
z��:33���2�Jh��?��|k����k8��p�ƾW/��&�t��~Q��ly�����&ꖵ��(���+����� :��0OydjK�	oBg�Ѐ��*M�����rr]�����y�*	B����牴&�ƌ�K�\�n�KYb!E�mk