XlxV64EB    3f83    10f0��,���"Ը1y���p��ox|�M��9��L��G��y��b5�h���/� k��&gw3D�<��r�Xbm �^�9� �A��E*��+v<��o�Y�w
F�j����D��K�kTP�"�"$\Y�����?`�NN�OU��S�"&7r���P�U�@-Ϣ
v?X��}f��+ĩ��F�Vؘ�VvM��ܖ����w�\H1������|
lã=-�4
����K��_s�i^>�C���B��mm:�	�m���o��]Z�EgT�8�"/�$�< �M���}O/x�p>����č\GR�E����bq��k��\��|���o���5z�XU0��x��=��U�b��"@V��/ߕ��d���O[����=4�
b��Ph�Ęr���ʒ	p�N��q�r9#���/�Z��7��8��B!+ôy����]]I�ad�v~�b(�걲��S�Ms��]c`�K?�{�~�984;s���C��[�=VI�Kv�EuB�n@�>�f-�^�(��>��5��D�e�D���������%��	�dv��]���9P�5g����<Z�H���ǚg�w;IN`�
5�Qu�:�xl�uxk�-��oO;H,v!�er9�a�}��3��G�����f��_z�� �㋠Sɰ���)����u�aj�ϯ�A~���\|Gi!�AЅ�&f-qVl K�\;��>y�G�3^u����6
>�.��5�c8���c	�!�@�w��?��u^1�C�ٹ��g
,�:�t�����Y\��i�W[/���;�l�m�2mN���W#�<�����`�]�:5�,ҜX�:HpW&����I�`�r�-_�����w�G��0�&�T�aP��3i��X� �R���:�KoZ�pY����e"H|�����>��-�oU��ALMDa>�-@p`���v�T�=ԹM�H� >gX�,����D����C��kC��,^rx��~D��xE\��x+��0��Q<M��ǯf��#q�|Jq��| �@���Of:I�� ͏t�����B"K��hI�"=�48'p7b�
r	&��ӧ�� K`b�E�:*x�Uo	~�4���ϑy5;�vV���L���ʞ�P)��� ie��D�x���5ڂ���V�b�#Iş��,K�|y$�|W}���t��a�`ݑ!�cn1Ƃ�J^�s�����E����.#`*L��oR�Ήa*��G}�뽒ܘN`ɴ0~�^�S&S�A[�W��،�������ă��k?m�<$W�����Ψ����W֭O4@/PX]�H5g��F�>�438�d��h�4�m1�-�,Q���]����v��MW�@�z9��#�$����v�뚓�����M�Ayأ�d��p߁���/Ƽ��xI�y��s-��q����@�����zi�H&Te
�=�2(r�nbe�p8�z�O_���t�	�`+E��ۋeH���Ak�u� ��3��ӫBƫܰiV���u�+�g@Cg��f^����d7�k�	əĪ #̄���c��@7��[?p��'� �f|7���1��!z�Y Az��ʣ2i�0z�K�9>�2����ٳ�w	�w��I��Вv�ti�>{T�̧��\f-��h���G��_Ogcz䗑A��#�0<�v�c�4�͇�3���pv�gS������/_��Y���Kb9���bRK%wѠ��pݓ
���.!��v%��������YW���n���ż!�+nE���/���MaI��&l��_.��j��* ;M�٫������v���FE���8P�}����۸Sz ��Ac6O��< ŋ۟��6�΃�����U�fx>(�SoC�?�@/֐��.5嚲>|�n����Xyť���=�법�Aqܹ;�K��n�֡�m5�_�=/�F`?�B?S-J��b�LK|Y�G�Oj��1wQ�kx�.��'�z4����^qf	�����d/w�	ѕ��Z>M��:=�F�^�.���{�M�}��YP���g��%ˌ�
�7#��'.*J�	���C{�ͱM���Y�R'6w��@��Ӓ_!�c���`�k�(Wo�q�ʷَ�	q+H�3��{�yS�������%p�l3Yzx&�Ju# ��a���pX����h`!n�+	�m1�$eyH��=��驊	m����lG�����0�Nd1�<fNaĞ��|����u���%E��(�I�N9�� ��}�l�U����_�¾_P��Ǵ�O���c��>B=��Q���KA��@ܺ�p;��N�`�F �]��i�6�c �D���5)*f'���
c��������iGU�k�<��Z�'�0dB8o��0���eح�S���y�0Un�4��<p���k+M���;ݢ�cP��tuI�gr� 	=�F�V�,1�`��խpX�EV���K�����$�ѐ%.i
���Lj��L��x��gQFu����B�D��k|F��#ۥ�N��w�W&l��� �������fF�c�>D~���#+P_� sM�)�D��ߛ}�u)�j[r��O����5L{��Z�T��*��ɜ�ʜ��������N����@�p��iO�w���8���j���y�7�1��W8���}�Վ��2�q�����r�2��
��h�0&��#�%RW����1w�g+�w��掜�F��Y���\��B��ٲi����>����R��Y���;���x�'�ȿg���k:�ga�߮��Ƿkؓ�"v,��u���(���,y���c����2U�f�!iip��˝ɥ5��4������d�)#��B�ó�6�ٽ���s��t������aƧ�A��pSti����y=$#\�m����ڼ���PUlC��e��(v+�|�N��w%}�x��DK Ps�"F\)�Y�X0;�Wգ�X���G��tYVfĽ��6�@�+Hk����������1���J���TD�]�|���1��g�i\5�"��r:4b0G1t~BNw������/�ya	��ǉ�Ħ�Z���S�4��AU�N���}�v\��{���BPg��jm<5j��r�M���W+˭gO(�8WX�u����Ϯ���ݵ��[���.SH�r� �2�]�U�!`i\+_}���+K%��3e(\GW8�Tgͪ�kA#Y4����Q���|9b�aD����'��Pn 9����Xʀ3S�LK�����T۽x���7Sw�F�X���(������W��&���[d8-p�M�jͮ^�.������`�<��Z΀u�c����Y	f�j���R�#���ol�~���M��у����31}mH2�-.�:���ޑbqK~:�y'qL�;I�|���+$��寈3c /�^�M�e�(����7Ke�x9Z�9��6��ގm��k��0�·|S{���;&鍕k�p����h�S�,<d�;���ci����pw=�Q,Ř�?�^�n	2�?����8{�Np�]]����Ux��� �OU|�`?�hW���S-�r�Vs"u����?��}���Ui�>���E	�u���}In@�{z���U��=��T�̌��TF��`�&}b��Π��#�ׇ��|�����	h�-����zWɤ���5��.bx c#HH!����b�ɳIA��!��u�7t�q�D����|H�� L�9�&�x��nqf/e�uh��d����c8��.:�:v��^Ĵh�LĀ
`yY�zò9�ߋ�?�#M�p�8�^�6���+��3�y�D��=)Wk W��*���֯M٭Q���t%��z?�4���=�_�g�(S�]�rI T�!~�V3��Z���n�K��'Oz�q�:y�\��.�����\���w��m�k�ͮ\��gw�J�dC���C�lt�����n�rȌ�R�P�䏡��¬v�#�����#�;�ݠ�#�i��ib�>#E`����e2j�L�G8K��iy����&:�
U���
m�.�����<�=IɅף	����p��6���Py�*G��������G���Pe�<�Yz�O��q��܂m�����'GAZm�\�>m�vD1G1#rjq���'~����z���CKfyD��H�Q֋�bKFV ���j���$���=�d3�M��\�gk~�+�:hv��C>i!]1�e�*'.g*c��,  ����ڒZH��Z䝰�(�o"�<�uiʘ�G�s�R˚�v5����ޔ�?(8�	�g ���G���c9Q�G