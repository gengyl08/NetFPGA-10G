XlxV64EB    20d7     b30k�s��̸I6��M|k��<�P�k�ܣ�Eޫ7�Ѥ�/o(][S����t�`��@����r�sƞ��N	W	YW/@[Fe��P'��f�[�VQ��G�_�B��5F�%�^k�n�C|����~#������!M)7�����N��¼E�&��ާ/��
�����O@n���8�Z�g�"��l�/����X��?�j�p�I����q�Q~}�ڃk�
{�)�����$��?�b{]�2x��� �f��>���8�~�~�SX�?����S�&72X(p%nrQ�{(�;&#Bo����e�D���7����(H�T�᭛��J?YH����( xͺ���»��TM�����
���0a:�h���+��D�Z����@���x��;H�`��-�r �8n2�*-��������qs���ڋ�ڿ*�Ī���W� ��iN����� ���)j˰�!W� �B	�b�=�[<˵���(�p�g��Q2p���d��� 9���TA��v{�Q\�B"^�������/`�{Aל
�9ylԅ̡x����'-rf�� ˎ����zӋ��^���LW�:���2��ܧw�:�� �W�!��l`��e���t�L<��Җ6��2���֙q|���><bc��R��Jg�&��-�⅒��Wqk��^?A�*\��<}��ڳyE~0ߒ5S� �3�#2��Vr=��H�Æ��^JP��ө �J����+�Q�A�掦wwߒ��id&��d,0�$i玖¨	j�<�3M�־���e�.���gK8����m_���~0[& �����]���܂ ~hK��L\��0���W8�J)�7�rv�8tJG��=��ۡl~�����2&���Jd=���]łZ��B�غ#�{�l�;ز3�Ԣ�\��c�a����̆ -Nx���A`yD&�m�|DSܲ���nuE�iv�J�u\ܵc���Ң9���"O�t�Q���\ͮy�8��Uw�����$Zi��A��=9��
��'���A?�emFk�Ue�(����Y����]�ʳ��V�6��D[�y/e��
K�0�a�]�0��F��
⫇���V����v-T��Yl1��`�X(�$���2�8�w��Ԝ�h����:A CnZI�>�����-�	��P�yߴ�$e�O�����Zd�Sw�᛭!E��qU=�G��*�F(ʇ�C�Wfؠ�N�Ĕpz5�.ޜ�[Wg���/kZa'����s���>ǃ�?b����� �{��4�lGlt�f��q��|Y�¦�b�\PW9s���oN����~��h���B��2���g�4l���U�M0_�}����k~RY��]1�(�Ѕ��)E�0���k�w	��������۳�PbpP�q�!iP-��H+�fT�;UF����ӆ{p�@A��x�;�%١�3��3T�I´��e���d&X���*.�f��K��+�?av���{CM򜹎��A���x�a�yl<�#f&��+����^1���\P4�d��"��t0����Ƞ���[*A[�k9�g�(3����j����X[���e�0�L���GD��_h2�n�u�-�9r,�kǕn����%��rm`��v0��QbY����{Eq#�ĉ$�;&� (^�|�B�,�7�����2����ӏdR!v�A��6N����k�,��f$ɝ��qD}����P8TL?�O/�v���_!:��"G��5�'����'D�u�I��Y����/�T��1w&S�����_D�iS'����Va\�K4�v)���i M���[9�5��^1ęy@j0՞ �z4gJL��)\�sv��w"%���;/�;�|�t���r�;��`�Z�����'G����v������d� �X�@�M�Z���Q(3�l���n�^u=N�=@LD�ԇ9�`��P�qlV5�F�fd��^����ެ�:��r9�e!# ��!(x���*^�(��(�s��1QFW��~��)u�a��7P�Y2d�Z�d��w�����}�L�\��L8�\Uѫ���k����[}4�E7~��ݒ�S��0R�kE{q�:-����D����v+ݿ��,���i5/��[!q��Q�����_��^q{�1c�!�z��:ѶD �/��!�{�@�[��<@ɥN�,�f�T��A\A�&�߄Ϗ�ϫMR��ٝ��� �Nb$�#�Q����)[��I�A���FJ}��6,M�5���mS�{��V�cC�SIT�����y�e�ix�3`�I��g�O]>�)d%;�ր�b{��`���`Q|�sQ��\�@^�KE��s6�TwB����H�X8��V�\�߶��;A�h���Ѿ"��<�*(�G�� Ѷ�5 ��m�=�]��v�U9G_�޶r��'��³F�����t.4�q��;��x�%���Qe�\���+�T�K�ͻ�(��T�ֶ��ң&�YcЁ!�$�O�֙80$����t�%�l )sq|N�q���{�g��a���&*D_W���~y��E��qx�DT\Wwc6�B�Oߌ����?����{�Z�&.�{�و�%�lq��s�̉��6$���N�eO�k�J�u;�gn^̢�b��uiJ�MV'�P:cy��-oW����ZO���Z�Z]��j�D�*��3l�^�/*�P��S�����K�F��}C>NK2j4Z7m��t�jj�Tc�A�S1)�x4r�F��VR�AA�K�J<�q�(�E�z ��)�~M�@z~��@q�zo6��>kH��[�A�XG㫥r�L��6��b0E��M�)E�ݾuG���O:�v}.��.��A6;��X]�h