XlxV64EB    3f12     fd0���&�M�_~�b��1 l�i��lx�����i��*��v����h�|D0s�Ns�¦9Yw�E����`n�Z`^=h�����9c����n�X� �y�n
�T�*Ȉ.�(j�e�߈�����˻e)��oB�)��Nr�loWpBPS*@*�.j�A�w޸�DR�}~_��$�N�no	#l�mݤ�L'��@Q���ޒ}��M�qO{h�u@��۫;�`�0����M_,��btN��)��Ź�����x�z��?�phu7)v||7W^%n&��.gu�6��-�.ñ^���|���bE��3*x����[:�Q��#��\'��`E�o9��mš0!i=)�Q� �@��ݳ
����15NN�!�)2�y��$�����YrI[���#��ȭQ���79��rU������D����i�
O���#�
��t#Gѹ/������C�{������W(y#a��1H����^ ��V�Q@������I"����MR�-ά�Go�J�x��yt��a�V`�����c�H~��2��J�/����g�l���Q'�?ǳ��$�o��]͔���Y��!���^��I���@�N���������OZ�M�K-%Cw�� D�/��6�ʈ/$5�����|�xgL}Be	h2��V�*�}��b�>���q� ̇���8MP��b��K�#�<����9!�c8��,����!�XF�i������ˋ���U�(X��~:m�����n�![��m6�84f ��e�Q�ݖ׹�0�eN�tLxE1y�T�jƧ���J5`F�<T5{��*>�;�!� 9q��6Xt��a�i��(�Ou���Xma�̏ş�?���a���l6��kȻ�q�$&�(�F��������wo�
�3ɕ�}~����Q�������Z�!��ZZ�@��u,;���~��^������Q�	�߅K���2���]��5 �>?��uT�?�zsM�VQ�7��*���ʺeތ�K�C�Q)>ݼv����G-���_�?;�	�?�B�q.��w����\�
G`�B6�VTS����΅� B_/:�c��Gυe�*{n�1�f�8x���hI4.qil�}E}{
8�G3x��J�C�g�7ɀH"��n:���.(C��Tl
�Ww0.����8��#������E!�Y��N�r`�־� Naa����Ew)q|�eNR�������d&Ňb"�u��g��#�͡M0D�Yu�`?�w~ݛL�u~+^,�"t�x�4_�:���ڼj��tM�q�;�	֚<��"�~��P��j�l��Fi���u��;�ՙa��c���-�5�`<1�S.���r!*x�u�U!�>҂��fն[<IPY�N~WO%��$A�L���kC����������f�Й�T���NZg[(@u
�"�J�CJ���ӽ�>�\�g� �Zq�E+f�b��i������9�\e���a}*�lĥ�Ԓg�"�=��U����&�RO;|��IݥÐ�惭`7_�����Y�쾸��A�,��]G4����]��a�3�B\�g1_���L���B�6ع�����ܞ�໑(ϼ�1�8�O�mzкv����v��wPp�.��'C�x*���!�-
M�T��*�C�V�g�i��h�w��z^e�q���6l��H@����ԩj�;}D�^+9��*��A�3��h𶆊�Y���7�"
mS���f	YP�E���F�引Dg`������~jv{#�0M<0�{;̴ɣ�@� ����)�SZ�I�-�z���^{��y٦�T۲�f�\�$�S��B��nǧuU.�Ϣe��`��E_r��YZ�q�p3�,���.�� �|�LGǕ0�;s��\�B�t-��,�<�^�̭��?����� ߕ�:�	s��.�_-��WD�0�@ѥM��]k�K9/�י�,lc���,�$�XMd	a�QI�2~B<�I;��g
Y	܏������,ߔ�D7R��[�$�^���Nj���\ȹW7P���;�L�M3��.�&Y E8��:_�z�U&&T���f�����G���9�%��T�<N��*�"���'XEA�*�$#]��~��!�$��=Ǩ�.4���0��/o)b %���X4�n�@P�ly�ܽ���UĒ0���^��Ų��cF�mf�៨��5��K;D����C�<�~J��<μ*E=�R2�_�V��#�5�&��ۿ�G�dA��a�S�\:u_!L�ܐ,YLZ�_�����J��q.�}c�r`8�U�Q_�GΓ��mɕ�H� lιBj�`K�i_�
�N��� ��43�0±�|%]��S Z��O׀�p;�|�'������Y����K�4�N�h�n'�'J2����e�R_��j���Zܢ�&4��:���gs��5�72n}&����nUq%����r�la�oPI�C8>C_ㆲ�p_y��L�;���b}���㵭J	��7��5Mce��Pl�E/.ǘv��K;I����[}e��a�Wcs��=ZW�g��r��95��e��H[p���3�f�����8gR��Eև�|c��g���
������0��G��&�\�y��ksMU������ġ�g� #f��-�5���M_��f<��WGĵ>xjr��a>�����*�g�-+�)�S���������<����G���A�	p���@s�W��a(&��+kF\J�|=
aF.�
^����N���Q�� ����RĊɊW��?'��<eŠ�����P�$p䐝��uq�m6��t���Ò̫�y�O��VO�EI��:��DX$J�<4�0��G7EX���!&�[������w������Ŝi��N�fv4a6��Y���eK*���/��Z��>>h�#@�8X�NZ+��\oe�W�2KX
�����g�QA��x
�{���$=,�Rע���*�u=$݉֩Z#��xF_RGjL��U�� �����VCc*|4���C=~�ؤ��;~;�9�@�G=h�޴�#���4���}F�~� ڽ����a����í��e�|����JS#U�ެ����-0N��W��e��AU���jsz ���*v�k�
H�ĕ�b`����"��?z����mY*=<v< 5Qv4ؙ���jT��\ }ԓ�b���H:�_[nVL�t9��7�du�.{��S����$�����p� �c�T�;��U=�HÃ�u��I�ƃȔ���#:V��h���|6��Yhɯ�Ʌ�=�3�Ak"�q�
%2���X\�����'�H�p&�H�q���Z���t�$�"�Ё�E������Xz�R���˻O3��ˣ_���rռ?_�`E"Q�)�O�oX7���w��{c���у������&���js��i�f��e����]�hy�k_��v��S��t퀟�"�mƫ����Y���S_Mv�EǸ5W�'����x}������Ui�F���z)�S����fN�KC ˨SWl�2�~h���V�F���N�l�^_㌑��ȫ,[n������@��S޷]j�5s�[�_��9�~U���#�Ԙ�_d��y��Y����0���B�orqA�'�%W؉���]�E���ЫhU]y�[�1x�T@���.���*�C݉.���&�gu�Z��~���}Ì{�cH�~�Qc�BD�!ʢ�b�%�cn��0�?�K�3�o}]Ҍ�H�q��f�ȟ`��7$�TI�][�F��l�ȫs\��b�M�eT8��5.!:�?W�=me�X"\�c�����̪��WI��E0̖륄"Q,ξ�[L�8m�0��`�$g�W�h7��sH��]ɩI��\j$Ӈ�P��������r~�zeH��ʩ�ü�r�	�9�G��!�0�|ڒ��5
��Y�,����]q=6
^x� ��\W��ؠ�.@�>C�R6���.���?]wbS25�{��(������t.r��À�=T0DKdl��z5��