XlxV64EB    2d33     a80	�
Q��!��� G#��c3�!�"�$��+dQ��]��{�s��2I��U�8��bo� ��t�GF*4/D_%��O�y�ΤLռ'�H⺭L���-���w-My�D�ޤے���}�нl-�3���������zz�p�L�-����*O�7�&�����!��?���9w�2Ib�y7Y�iU�x\���]����V37r��X���kPrt��B�J��P�<<x�`Ǚ9�Ƶ�'��#�$��:=|k��E���۸�,�*�cd�.|��m�!�u�� h
\��*`1P��5�;%8@/�kHEbmr�#3y�p�9�ɮ�4�3��$�}�"( ��c�&5w���?%u�S�X�Ed�̿������7KY����Wnz-��Q]X��2�vIkjU�]��C��|���1�P�d�T����6[��>q�+_��_0P(���Oej�(v���VZ�"4�n0t�<-���WC[Ր�M��~ ��J��C�ʨih @5���i~�ň���y�@����L��2�Z���`(j������˹RI*�-�R+�j�u^/��4�e��o�<�QLJ���.�,�TŅ�n�d>��U]�h�����D����4{��2P���u�6�K;�̰�qeN���O�ُ�Mqi��;�ڃ��L���S��������0&��x����!Y��7��+~[�:�[���!�2Qkw\�ص�qg��OK��y�k����p�Z;U0͛Z�bo�Mp�wZ�8�wۯ�e�XZa-d����}EPX�3r@�MClz���cY��^o��zL�SN����j����6 �W�/X�:�h|�Nroag�/p��5�lf���EDو.�8���ȟ�m�0:����A�Ҝ�'�`����ܻA��l���}xPL���@�jf����:�I(Y����r���c��r+Q�~C릈�2e�P�FT�=�B�H���L��)��zՓNAA��eX~����d�p����t=���q0*F��m�X0�z~��0�el/K�'D��Z���T�������w�Whb$od%����	�:E����+%G���kS4y����|̅��&��nB��
Ԏ�Vy��ܯ�Đ�(>9�V��sA!�1�Y���0Gu��Bk:�ا��`��u�Ay�\Cl�5�X��P�9��}��tJ{�n3���~��l�RZ����F�2G����n�;u��) "{o����=F�<U�����4=�B����_O'p�;ñ�X�n����eS��+�yC����¬��\�9�J*����A�,B�Y>�A�,h.;�@�|o�נ����++��
�D:��K2��&T�(d���Rns(`p4�kph�(_�\�ŽI�2�<ŀu(���?[��,��+�(��7�I�0�����s�����tI;�zti��䨒}��SMjA6)�E�\�f�����Ќ��0�m�7i�b��E9�>E���	f2~�a��x2�/Q,�K�o����wzqH����?
;��@fG�� :�ę�}�`~t�����Jr�U/����g[��9�T
�<�F������O�jr�:2&��g�_3?��R��"�GǷ�t>8*��� �F;����ڊџ�L���;'q�æb��:�Va؞�t�n����^�a4�1�Gʗ4�=r\&�J�MVɱ�@��>�m�p���|�"�b��`+��W�d�H�8��E��_]���S8�T`s~�w�3�(M��h/��������ۼ��U �)e�wT��m˯�L@jb�A������d��,z<�5uW��ɹ
I��*O����F��ȅZ�
_>��3�����Z�"Z� ���pv'~S�/�[�H�W&\WQk[�P��w�)�RB�xls�����5� �+���0�m�V�G��ţ�b?Ϥ+���Aδ�3�!�W}4:3��7n0��Q��������O�fV�_.��M��VU;��w6��]� ($�)�þ���������s����ȥ�0V�XD��z�Ћ�1(7V�H>�i>s�i)E�$�I�H�_`�?3�1]�e$^'isR.fr�šA7+%Ϣ��r���]�n�3ѹb�oZ2��|��̧��HR�)�X�D����6��T�ۏ�/�m��"HI���X���q����b)e��p/f��U�$�܊ק�7�v�*XCDh� μB#\+�?�'d����덂�AoFY��TX{��p(��t�7J�3zj��l�D|����Η@���B1,������Y�{� �Đ2s��] j�^�F�����I'<�������~�,�q?`V���ZK;$�o�E����k���q��7��u�+��s��������t/1�sq���)�(���!맻��R^��V�ƺ~�7"���.p�I�� '��y�l����R�����o�@0���-\���t0-�[0Ev{�䐊?�9�*�i*>���2g�!+x�� �a��ϐ&��!��w��H8�%ia�hD����p^c����~��8LDbhE�����w�F��y� �1S-3A�P.䳷:mER�R��bW8� l�|�pJ�å�őZ���b��弶�#�}�e�ه�;����yg��]������V>I��i1��`�4ɢ��l�s;��p