XlxV64EB    40f8     dc0m$H1����4�DSAq̩����W4��$	��c>&���j݊���̪�u�6�}l&��t9$4�'0uf����`�&|k��^C�L�1pND�ɫ��X�d��nO�v�%�}�Tp�Ү�Hj8���(M��������t}���Զ��rZ����]�!ٳ�����3���l,2���2����ԀA��$%�Y�а�.���}��� �����2c�϶��W�Z�|c����<Z��SN���Nq�XT\"h	��:ɲCR�Z)�K^6З;�Rz=�Q��x��
����J��dk`cU�ɂGV���W��D ����GĆ3�B���A�.�$+=WI���A�y�)`A���G�L;G����M�����Co��#.�!�R�d\�C�{!AŴn�̌����������M����G���.�c�w�m�Nї%3ss`��EJ��fWy�\����S�9��0�t�M9�݂6y��.$g(^I�V61�2��%�cn*n��2
������w��xb6F�|"��W[��a��_탖���ẻ���~��#�U�(� �*&����'��s�ն��Е&`�mt��(S�F4Y��j�F�EY�n��ˋlJƆn0@��[�(��1`��~���@�ο�<����ș��Q/J���}V8z���$��;}PA���^�θ9*�/֬n	Yٚ ��� X�(-�/�O��)1�Dd}��q=VU����v�x�r�&�Z��J|O����!�������#DRw������������wlW�<�w�9��3}�G���'!��ڰ�G�E#$��1��K��Ud��|�����U%m��D���	w;;6��]��� >�j/�,�oTg���^W�J��ɡ;����I
��c�sJ�쿂���S�M�R�4��^ �-�g	ʿW�Ypnv�>m�ϛ�4�`ɬb�5�/�,�e`��Yj�=�m���K�(1���{z|jv�RIZ�I��X�Ҿ�sp�O���1��� ��<W�u�!�<�P���`��}\���L��X�b/in�NB�6�R�Z�O������
5�L'�v.*��/�sѮ�!�����KiK�)u��I�����tI�;�ɧe�=T���a�H�0��n 2#�w���6�|���0���E~T�H��f����dZp�U#X��\=� ���v I����|H�C4�`��C#	}��=�:ϧq�A��0�a�4�u/k��o�0�c\%� ���C�%��mS}��M�E7� �����Q���+�b�oD���y�*��ܴq�v���=���@aC]Z�Y�Ծh�F[0��sOI��� ��iڂ��d�!*����O�<��NP��[�hҞ)�R��y�V��*8
����/�M�f��H�	<o�#�lȊ�<^��!��T����O�����3@0��g�串G?6����+��x�8�H%@��@�B3h���d:$�X�Z�g�+�e�.Z;�U��D�Xv(��һBU(�������.��ڔN�Ϊ�h�Bj�Y���>��1�O�~{lJ����(�i�txv;ۮTTFQ�'G����22u썱/��wpe���� �)oh�l�i�YcYں���ʸ�Zd/����쒮Z�=Օ�xGދq�޾iP�*�q��e$�MS�yG�j�r}sՑcX�Ȳ52i�v��<�)rX�]��G\�p� 1ɨ&�X]T�&�ίD���h�/+�����0h^w��Mj��+�#1�qX�p�;�1�/�'���kh�we0 ���+"���(?�$�೔�w���v��V}�ϱ�_���@�oj�����eø&���<I9�=v��OTj��q��?:)�Z-e\n�4�\�}�k	�#��3��t���%��oQMuUZ��:kZ�`�B'�ӆAϓV��,>e$�j�ώ�?��m!�|^�>���k���8�p�àP��5"���
;I���f�9n)��}��1Z{�n���Nh=��qfh�U�B_;cjb�xa_�PT�2ﲈ�ܻ��������;�y� ���؝��*rq0ci�ĩcZ�+9<A?��h)[Z��x��}��T0��b$��
x��t=�c�a�?�{�����Ԏ}���P��|p:Y�+?5��H� Dof��H�v�Ș�cB�*a�"������y�ӏ�܏b
51Q%ON�;�����x6y"�<x����C��������ڜ��0#�j��y����2��	����^߷�~�������3%�)a��O�� !��٭J��X�f!j����W�k!����~�hf�Нqi|��?��dҧ��h4O���`a�D���s����Q�*���X�)���d���۟M�ty��(3���b��-���+�H�7G����	4.�ӶD��D��׍ �(��}�� ޮӉ�~�\7��]7J~�|V���$%����RHX}E���B{�����QE�I���?�Ւ�'�<��������T�}����W$�Bg���6�]�p&%�K`u�/Y�L ��Ԗ�Gw��R���M[K�����~<	�,�<('�w=�#{�:i��B�n@:׆���h��NDN�`4�xu��F��Gs�\H�񶊍�N�t��V�J�ѿ��ˆ���T8J�aI�����G�y����~�g��yʠ�  ���[k���V1����F�S�]�s%�[��;A6ka��n��T+��|�|�A�M�6<�O7ҥ�����I�n�7 ���tT [�5��$�e���K��,��KP��?:Ԩ��S�|�GT;�oF�x�N����I�RSL>R��R�J��5�̲h�&wT��\�3~�f�د'�^؋	�U��cw��D�;�iD�>-��]��*W. X�����!AC�BNF�[Fj	��߄uc�ܔ�k:;���3*�#��|�� ����)��@�=���z�C9�*L��5��!&VArh��bT���~����Ռ�|�S#s�
~�2ۨ�����:a�׳ͬ��R�L!נ�&tJ軫�Q������b�G�!a�s���o����OC�!�'�y�O����xT�?WX�s&B�����ę� �����7� ��~j��1� �@~���QN���ⰞK"~�N�v��a���vf����;�n����y���Q��R�9��Z�Tn���HM��E�cl#9e{ ����D��Ki��0e[E�͖'i+�H���9f��
���R��Q��|:�9H����=�p�4x�FCNU��L�*)r$�lf��1bl�H�W[=�Z�o�KqL&�ܡ��ub�]�/{����l�r_��Ӌ�r:6��$�k�k�D�M�z�'Pf�W�bp����9�^amv�ӺZ1����u8�n��O�Ǐ�k�gi��g��%���F�x8�bp��G�