XlxV64EB    153c     7f0O2k�[���r�%i'�!�^�Ŗyg���z皔��huX�̔�l�gTDX���ږQ規��� h���<@9H���;2q|&R4��C��t���g� �]`y�0n��f�\�z�2��9���|a� ���o���K�n�e�=���O���c����bT+�6�U��k���K_�l�q�2o��+�2�z������`�HT�g?���ׄ�:��,����"i�.��{!�4��t��3�����zF�˲�)f��I�n�w���K�6�́G��m�bzAu;�W�w��1�N�=��	�v>��Mz������5�`H^Yݳ��EB�i(�eX���c���Gu��H�b���4 b!�x����k��4�d�5D}F��/c3�fkn������nzm�x�@=�(d�"
ػ��Y�#@�4/I��F{�w�JB�n)��J���U6�Fd�K!�r�{�}�Q���:���=��7����C �GP�L1bc���%u<M\$��>;t�����m�4M��C�J��S;�]$��B6�'�����^������\�!�d�o��+�e�D9i��r�v�L������図~wl^�*S�r�l�
A��Ls��5$�"��v�Ga��[..���,�����w)z���*T"�tT%zgQ]+�c�ݴjY3m;�����EA�+�(ATPx��Yx�w� �'/h��P�'�"�VFX�����Qq���x��������,��,��F��N��7��%2}��Il�H��� �(Ӄ����ʸl&K���~ua�a�yy����Y�-��pI�ͽWkOms����[�X9}�����x�@M����G�rt���*�bn��DCk�J�1��V�{cl�i=�6���Z[��W���8i�����L��l����D����;�2T���T��i����t�۞䊹S3�OO4�h��2bw�܀���8u�>��m6�^OR}������Kú	��GоپćX�*�h*6�����Eކ���G�֕hl�y\��d��*c�c��~��DY�hA�"O���'QW!C�K֣�C�S�R=+ړ����L�lv�#	5��ߗS)j�>���͙��ˤ0g`���N��7��$�W�1�z���R�J���`A����Sv
!XyU�D�*�W\v��p�pphf��v��l~�>�54Y�`R1`��R�x�w����4��B=�l��g���Mޯ=Z��c�p��
�s[�L�V[e��"t��W�$��&z������hjrB�l0)�?��q�h���'��~�A�ܫĶ�Ң]��h�:���0�_�6tFBM(��~.0'9vl�͋�����$�H�N�%�p�@WM���˨"`�V��RSuB�"��Hz�Ĕ+����A�H�LB���K�w+`����.e:8�s�5�ͪ��ǝ`��{���Jŷ0$o�qz$,)�!��s� }������|tS�j<K]���u�<VVO��p
#<�_�'d�´�;��g5�W����f-�^C���D52�K8��cyfȩLk�2	>T@s��/bu��G�ype�:�*��N���8t�>��5���(\���~p�\ک<��Ą�����<�>��i���x��պ�������Ea���/�M}���56��E '�;ϳ᜿51� t���6j�+@��c_b��y���Z�M"�b�����;0�w lx���E���������v; ��Hw��E'��^{��Y�a������X����J{<�YI£ik�/D�o�|��d��������3֏�5��a��_�}J����}L$,��K�i���"���6�����%Gj9�]q�5�����,�j8�z�K��GZEw��p>�Ly�$�\#@:��꓋��Wp4�rs�Jƍl&o$�q�3/��t��3[�6㮒�44儬��K	�pEg�4�	E�)!(U9Wkg�5M�
�u88)�y