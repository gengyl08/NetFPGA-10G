XlxV64EB    2c29     cc0��.F������1J2MZd�7�J?�/z@�zIVY�ʡ���RH\�����:,ޑW)wY�l9:�X�#�[X�,�U������ג+�LR$�A�0�o��q"G���
���W���=�}����M�Y�<�p��|�).��Z=~�d�e���tΊfwQ�a/�@!Q��\���z9̬�i�㗟˦�͊�kx�aK�oDӗSRCJ����-��ut�s�O>-�2{��p�OG<��.�5�r�@b��t��jwLz�`� gB�=��>��i�����y�x����F*|�p��o+�����@�P���*o
��0v:_��/�2��Է �BN��&�#ӳ� bs�{me����oj/�έܢ���n8�Cd�����25�X0���A��uv�.U��A['O�i�/��m3����H����/K��ø�a)H�a6�gC��0�Q��x�誨4;���r({�u|��K���Ѯ�QJ<|5����g�#e{�/��.����~�O�F���3�iڂN)v����ɴ��YV�����I��46\Ը�U9Օ�W�k��x�Q8ˇ-xO$]��,����V�Qt����V)F�u�B��Ћ�!��7ǡ?t[!K,p����i9�	W��+_���˄�d454M!"��:4r_J�F�S���F�y[C@��*�{�"����ZRi������Dt,�'��`s��wy4�W����nC�K���/7쭟�%:�ԇ�O��yZo@��2�,^��
�����)���D�l�)'`w*���H���hNR2$��jd���l|"
.Ӂ<����[5�Q3��c����RϘ�E�D��:���bH��A��R����C.9�BJ�}�[��۱�#%]��m���%Z����j�P��FJd����1{.�҆c�TZ��Zɿ��R���.גt�����)E�?W�n��<��C���O-��-л�[���k�G)�����7u�����С(W�X������O[nF¥!�K����
�ts��7�=��ʈI�7�`�_�X�ywD��d�V�u!d_��0Π@�F��{�Q�D:��FF�eT�bȅ)Nh�(��6�｠���	)8F�����f<=�#�Ty��G�"#oB���Q����V3u1��!,���Ӓ�
)L�ѐ���l\6���G��H��\"㌓��̗'d%��|��g���v��H �F��
�����|-Vf���ݗa�2,��ǟX���!n E,�l"��A� ����;O�W2r��\'��g��̛Laх��j�P�	h�59o0
8.�0�Cp���%5^��k:���K+�thޜ��P�ݙ�6�����|��Z;��������r���D�
��� d������!֜D���ʥW���a�|��(K/ONowS�
!�e��4'sX��"���tR�x>�8D���.5Bs����5���kn�A#
E�_a�\hL*��@��`4�8�\\ĕ��q/C���^��E�x7;�"�.�Δni=T�,l��G�~=qBA����08�Ms��Ta�Q�1_��VU:�-O3a��kC.��^*J�!���ZZ�ۯ9���|�3ȉ���2R��FU��5�bV��a��Ja:w��&��^qΫ��RP8඘Oj�yҞ�Q;ěğH�3|Zߍ)���TYH#�/)"�'[L
���|OT�F�1I����K
)�M�+�J�&��]��$\?��dJ����}m8�|��6��Ua�YY �D]���6���&S%.Q� ����&/�
!�NR]����-��J���7d��._>��ә-_/DVo��uW?4�Є���W��<��av��T�X��eY80wP	~ �q�����������uj֪T�_!�����r
c�Y'��O���/� L�:��'~�jQ$ە�h��ӷ�b��y8�5�	fK��܉�1�����91�q3�Xă ����}w����E�	��a�G5�5�t�ڔX@M�C`6�Ѓ�k�`����Z�c���C���.A�$��K���˜���Ď�[NN�K�{=k{��S�2�s�Yo2SQ�6l &�<3��Npy/�:�Y�Q !u%�	(
�=��S|r!�9@i!����kƋ�<Ɛ�qk3����hI+���@���8+~{�ܦ4��;�`Y�5���s��p��`�l<lr�;�}�����z'�'��^v���Σ�gۻ���8����T��@�S���x��������\�\�tP�+���ff��]�{��I31�C��v�n�͆x_\�F��&��c��y���C���{��8�K��g�8�^�´����}C>P�am#6@=�2!�;>2c�vp�#B��>ߓ��"��������Ш���<z� 5㕇�h~��O
�B[�����d��p�<�K"S��I�r2�#�� l�7Қ[,���X�ey�{,ԇ�C�	����8�o���U�|��������B>��F�(�4�x�=`���QP�ќux_��%[��u���h�<�:��=���d��Cw�~�}5�p�Ƶ�[��*\#�`>�.�~�9����-�1��d6�`,X}@��f���hq��R���� �j7�#\f=�Z��{�-U����aJ=�jYv��ڥ�wM�z�<��:��ld��+�>��
���Z&��D��(k�'���C�g�1#%��i�S�e��r��zdM*�$)8��hf���|���k��O;�z).nD0ֶ�p���y眼4X��)��+-}b$��G�R?�����ҐV�3��d���Mn����B};��x�M��"�r/��껺w}&Y���jH��������ż��F�F��V �}o��鏤.O�ϟ��:��(�hyw���7�߬Q��ڿhRY;Q�xu4�p+%_��3X/ ��8�
9�3e�H4*������B�� ��0���������1����V1%ND5}p9�y���FR;��o۽wI�� N��N���/��^�BK���3x
Js;HF�^����@ŎO�"킻Ù5�~��)�{9�3��@�!�+��
��D�*�r�����1�-/�֜�˙ ��U����(Q�frG ��Q	�.�̺���n�
s#Q���H�/�B�����p>ь|�~aJ4�%��m��;�:��� ��%��Zݢ�-I��M��Z��;�wA
�
'>oC