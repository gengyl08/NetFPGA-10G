XlxV64EB    1e53     a80����ם���\��=��e����V���2�:l�3(��m�i��\/��-V���N������%]>�>���v7\@���o�Q޴@�8�]���g��Q�W�u�jӺp��%� ��>
Y�_H�>ű�}I�s�Ħ��1���,h��v�����&�Ď�Um[��f3���<�L�-�)Kf�L�Ţ�Q	�t��x�'m�y̚I����?&(_T��zۊw�ɚ�Mp��+�s��Me�瘻�,��r���	N�6)����wk�sذ'q��rʏE5ڼ	�G�tҫU�%` (�<N���E��&�D��3�"c�z�6ز��G��H5�T�� &�LY���J&t3C��O�3���.������S��W����v;޶�,���E�1��Y�,�~/�j�(3�Ԣ�!b�5��ls������ot�V,j���8�D��sya�r�r�y+s3#>7��k���w�>���d�f�.s���A����p�������mU��x�M�m���6q-��n8�:_���&NQ(_=7%�S�TF�"��t�����cR�NUS��F�8��Y<q}��i����Y��s��٣�'WP�P#��i�7]�P_g
�-&�]\�2=�o=�o�`l�Ң4<�������kv�Ay����n��e� �΋�*�:��Н����m�0����|�X�Nb�Ks�nIw��<&k3&��R=G�6�I���Q2`����C�sU'0��Xi��>��#���y(P�,�5�iJ�b�!�4C�@}K`�|��6�F�=�%�}�{�	��b$���nc����oȗM�H�*���y��*s��-9�u�je����|�dns�K��,+�g�sK��>���Qnك11o�r�����s7.!���nL���	p>�������3���Pܻ��6�Nyy���Uv��W@�H���©~�Q��z��c�a�"��B5~�=��eЯ�)bMZ)�>k�K��^�P�b���^���6�g�%@�ھ�at􅱙�tT|�_�h�i[%b�`��~s1=V�'�ȩϭ, ����Sb���%���(��?M��puI��O�'�U/8Arkaft��\�n�U(?�맶B���.�;�4Ϋ�w��~y�� ָ���	(W��|����_���U
0Js���E$� �$Hw�h�$ϫ��8u0� E�z����S͗��49����h�����p6�.��R`A�J���;�U��B�������+DШ��j��G����[�r`�����[�d,l��X�f�AB=������NB5b���!�L�Pr/�pzl\\����j�S�O63���g���Cj>f���F�u��x��m�&�nq1(6b�\���<��qLA���2��A������UN��5t�Ǵ�)<a�~ޫ�ъ�����jp#-�p7.��-v���!�����ZOE��uU�KE(�ص? a��3!�G�̥��V�9n+�����5\��Y��'���F>@6<%y�e&�nϹ:&��<'_�_��e���M��k!q���so���0����!-E({�Y�}Bϖ,�~=��@E�3�t(�ܭC��1�	�?:\���;i-27�o/hr��'[��B��ݾ⤾�&K��h6����ܧEz�QM/���±c�� l����d0_��ScTi��Q������ﶒ`ܔ����N�d
b< �?rw�}6<���Z0B�#k��3Zж�����f��o2���

�n�?H��`��YQg�[ۻC���*B<�J9���<�j 
�^5�jx<o�7�<=S���)]ؖ���|cʊ�Y�K�>X��Q��X5��("�-/�5�	�G��O&��9u�Sd�H�Q|ws"�F�suZ��������o�M�̥�*����.(7��8�t5>|����/x�?,qֹ�q��b�7˶�$@�u����=��5��H���L������g.q�$�Ұ{���Ol�����e�����7)Ɲ%0G��*���?��P��Pc;Qe_�K����+�Վ;;7H7gk�#��9ޓo �Z@�yU=B yȼ!�BCݿC���]�|���*a��q5)K��/�~�_aA���ѱ��;*��{4�m~_p��b܎��(e�����!<Q���NWR�C� ~�º���z�q�s]#ed�M�F��є��+�
�a���2A}�]K~AEb���[R�N���~��1hɛJ�KTu���.��}
`��5��(���ߴ���9IȐ��=�ƶ7y\h#8�l����7�9�緽N^�eo�@h
Q�5��������{�����pߎ�������@�
^n�S?� Q�ɴ{���j��MX��wl>6��ؿU�x��NjtO8�l0�˵�G0IQ�ƹK:G�q�����	�� ��ly����Ӓ
������h9��ވVX'BsG�H�.�Gr@���QE�(1�B�&���q<DlƦ�]�L�8�m�D�U
rrG6S.���p-�(�D�u�웽�d�+�\�@���٨h#Sy�?f�HN�F����T`�m(�����char�7�
�y�~WX�B�Yh��m��#�7o�o�O��'�}�}�OBܶf�Y
��`g$���.S��