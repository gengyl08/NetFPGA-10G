XlxV64EB    5cf7    10c0��kӚ���}�u�XF��ӿ4)qpWHQi�
�M�"�q=�h;Uç\_���وm�4V�� ս�j�pYC^�}\A�I�A/�[]V̳x��5���i�9F��ѠQ`������P��%Q>� �6>��#�Iү�V�6�)�$������\�J6�`�h���Oc��L�#b������
3�2N�#j-�Alev��Jy��+׫8g��KA��ƶ3����%C�x̗����_�0?���1�s6tc!��]��M��T���=�W;'4E���Azw�F��|�kA6�[���کP�}�3H,��+��^@�rb�.�7�l�͌1l>�5�W��Z�fU�]�WY,��ǛQ�	R<��	�M�D����dc���\��T���,2gXJ�p)�KG��I�������O�W����=0PI9<Q5�$n轨e0>Q�S%����_sM��^�@30�E��4Ew0X:�<�jHmC?X9Е�NF�n�#�6J�A�f��3-i���S<�7:�^�'=L� j�k�M���2�Ew�p��u��8-!�T N�zI],� f��5r�FN6�d{�ν��Ȅ��e�OICN��U��Ň&kď���J����^���DX��j�3���ʱg68Ɲ��{���gГ��zJ��]�Q�| O�h��K9X��V,�p�c�K`��e�u��|��/n�Y�[�'�EA�/+�?�gd	�%��٫D�A�����Y�~�(����E�����N���'��6�]"�o� �pѼr0wz���Q�+��XƞHzG �C/zdy����T6�=hͬ^8iZo�
 B�;R@�2h��7�ʫÛ��-G9�'�˼�k�`?O��3^��S��=�B��:�%貺�b"��
P� �Zo�����b��yN*�gu��(�T��ۡ~F��О��M����0/&�£�'i�����ղL-�Ă�$#�N�Zс�P��[�I��蛈�4`�*�0ฏ8�`�W�i;�	3�h�u@'�C+�;xo��‐(���H	f���f��Zt�����҅*$����!��2̭��]	y(_�r�z�e����j��� ��C&�}�������B0��ü��2���L!�ӄ�Ј�(C�%<�)����i���-M-w�;���9h�.�{��;�Y�"��ż�]�kA��N7�0&�x�`򝼈*��iZ�**}�� <ߑpa�q��z%>���2h�^0H�^�G3���`�j��PlsZ�9iQ:���#��ZR��H��9�Ȣ�C/�g�ɖH5�vрQ�jE�!�����f,>�����Ԍ����)�Bݶ�>Q��ׯ>D���BEz�C,���������8��dzNɩ�5�6)�2g)�=�$�t������y�'��׭,�6�˩\�6,M|gd�)�56�`K�k��4t�TL���d?�X�-I��������M��B{�����9[�|p*ؒ����\�Af�k�x�bS�Y�v=������H�NR�T0�HH�p�Q.e�V�]d�V��f��yK����8N�%:b��y~!_4�%9C��XB/�۪���r,�ޒ�,��R)s��c{��mL�\C���K��	\6i}���f]����8dt h����R:��	��^l�����Z[����h˝Cz��&��׌��!�qL�k�9&_��`uo����"fڋ�o♌�P��9��u����� ������yd7�v{ŉ-72J�	/��@�p���I��&=����<U����vA%���g��?��dć0B����i�Z��W�}�IGoݍ	����C<+v��{R �bMk""RۖAG����L�״@/1��L>�Mʊ��A�B��c7��POeY��iS��¡F�%_��o��[g|�d������	�+��<԰������q�,�ӻ�n�xW�,�Kw�-�e��)��WTGM?3nq���*�l�R!�*<�w<>�@SӮ��ڋ|��!�Y��\G�Lu�)G�d�t7%*J��I�OC�oF�Jr��1������ġ�?X��������|�_ ]�g����d|?�44N_����@�������>���M-&��2|��у>�$OC���;c��;��j<��pL'���N�6mdi��ͭ-��PNP�Wd�)�|�� ~;a�)��bK�2��h_�F'تbAu�{��� ���"{@,���ǡ1f��k�ƛ���.�\
���D'I��Ő�����2|�Lp�/n<ȼ��+� ��%q.�{\m�Y_��w�f�co�w�V�a��L���I���롔�(�k�cUi&Ǎ����������ofv��6�������%3J�Y}C�Lm�L���*̦aQ�Dy��b�K�vpۛ�<���c�W�g�p
���8k
J9����9֍�`O>(&�	s	2_�X�!��1b�:P� �{��.�Q�U�9��r����	ѓ�6�����"sh	�����=������Xxa�{�z��������iҽ�q�֧��x.ϙ�V�A���й����zЅ����e��[-A���q���>��Q=L����X>ħ��Ӵ;W��5a����g���j�]�E�VI+T<c�	�w���qnA�K��33�}�4|�X�{F1��(w/�mr�)n�G���/���n4_�Rb�zrx���H��P{��0~���������O����N��>D���(�6_�Ne�5~�a������/�Ƅ	��?��^l!U�X�,"��9ݛzᱍy�]����BL[H��2Z`�U;�Apڒq�����������wr{�	X�l�R�*R��18xkz���INә�e9̲�+X�/O�
ݞ7��YFv�K��v�fo+�f�!e�?�
:��G,�n�T��=Kqu	��w:,X�y���IH�=��%Y��K�{�Ƴ�Dv��(X*��#��F䖉G.>(%܆���7�M�8B�ۧ&��p�@d�b,���&cor���J��]1g~������&� �
�Qnҍ����4�<�l��D`v �����9��$4.�\�8؉�����5v��CW�򸬙�0����SASË6��A�T:f~J��tœ XA&����ȥ�d���=[����Y���(�P���\�w:�)����$��q��l���	Y���X0K�4�9_���w����_ȁ����/�!�m���|�6�]���	�V��#�'z�B����œ2�������t(Z]%����V]�o@��ܱ�]�F�g��\�3S	���xq����Ň*rg�U�_k;J�wH�y=^�����MREf��2"s�uk?q)���nH�sy�<SP����Z �@��'dL�&֫��_�54����a���<D�z"^X���fR��8ț_i/E�\�:�_�kd���vRJ���ꨳ�3���+"}U����OK�u�"ò�"�LV���Z�k�&��D����.q��d3�;C�,ʜ7�\���6�#;4�.������Y �Ϻ���BnC@Ǩo�{ÂA�?jI�-��l�w�#iw<J33�ww���8�D�ӣ �Ӌ;��q��	��Dj��L�������np�ݰ�r_U�ܐc��lz�2��E|��V�	؃���/���'� ~b-W^�����#��I���|{�1 �|�h�_�*��F ��-��GL���<��TP��_��=��	у,���3'Q?�Ir;2^�p(E`�J���V4�Q�֓� N�3�P9[K?����������|��}�[sn�6���=�H��%w�87)����|��,mW��T��@��1�k:���b&��a�S���T���  \��&�	h�h���!�bg��P�?�7��^5Ҝ�Qs�&Cb�3�*� 
k�I3�z�f&�۳���h{ew���Ts�=�j@�S9���c�]���0ĕ���{���h7~ֈ
��[�d��F��(I����/���Q �^�7����������;�I�x5��^�E���'F�d��t��G���ڨ�2>�ͳgwG�v'Y�6ة<�ВW�y�)�P�{,�6����s~
���(4y����&@\,yGίV�ms�3�4r7G�\��z*K����+�/��Gi��hJ�|^_�E2X�P��^}_9��	���� yD�7��$�I�L+G�V��A�Y.�
�G	����pf*�*/�[\����Y���