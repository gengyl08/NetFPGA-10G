XlxV64EB    56d8    13d0������шm��񹧘1� <��|�]�C��j�3�3���κ>%��7��˪4�nu3/s�w�ߊ�}��%RӚ�����0{���4��E��+� ;z����PaH\5�̶_AKiǠA	Xnn�L�:�K+���.ewb|��q�I�D����fz_A�ي.�����b��l��f��8CT��sA�@,�-e�{3��PEC��k��4��.V���z�n�ۘ���D���^�3o���n�q�7�7��5�{ $6Ѕ�ƴ��a���^�5��0S@K�d��ݔ!�����t�{Z��3 �jD��(���t��S�︃(q��'54�+0H�)�,@�Z]�J����a���zy��j����7dK��GC��丑4��h_f�
���'��w���|@�[Ɏ} ��';Q�,�t�	9jҫjˉ�D*������Ǹ������"|Sw��?���qhh�m�X�D��f��Cu���?�����(Wlx=\���$�A�~7�Pn�}:�"�Kb!5�k�+�[n?$9&t�߻LM@��Nu�ū���xzl���礘Ӓ�������jC� v_����3������f��7���~!2<F_2���f飞�܂X+]$j��EINas�Gu/Uꇅ�S�R��x�>�Y�0��_]=K����o�pPWK�r�z��F�ʠ�Q�8e���:vm��o�P�:Ho��b 8��#��[��I~�a;
�l�a6=�RP��#�zlH�bV�r$��/�PQ�c�Kٵˋ	_�/�չ;�F�vU�[j,b��Z���_��
�˃�Q�TdrT����i8�x/~-��^Dx2_�(���VyH��F1 9l�����a��ܵ�U�[�;�
�	����r)���X��k���*���}��v��j�r��S�������k޴��b��X�ݤ ({Z��B����;���%1�����1�
�S���	l��Ч־@LK����1M�0�C��Z��ɸ+8=+r�y�޶*p�y��z b����8�SWkUm3�!·��jMPS��'�� qX?M�;��3XU��3U2��79�"U���=�sɡ�\]�S�ϭ�A���t�[�{��cEW�uD2o�	Ym��=m��%U)'�IPr0Jb��QL�%���,칕����H��u���K�b��Ey���y����[AE�d��� !��=Be}��5�[G��ed�"#��o;6s��cm���r��L����Á��
��G��D�3R pq���$:�3��4(idQNS�4��P�`E�2r,G��e����I"���s�	^gQ.m��a���m���}��E�Q����
�1��ru�$b�Ý��7�)4yĘC��=��K�ٓ�G�v���"B���W"O' b�"�ɐ��.�5���`~��ê��]�J��5/z�G�rs9�ɦ� Fq�EK��j�̌d_Oә� �[p���Q�uf�~��3*'?����f�Re�\lf���N�	k�/��;D[�u:9Zz�f��8�H�2D������jP�7~}U�%4ճ2�� Y��,wC�
��G�w��qs�M�i����6�L�W�+ӒW�T����1
,Bh�/�"_�a?��P� jӦ�lfgv�ݝ�ƿ}��#?=�p�ԛ|��A����\b�J�!
�
8}�')���Y���{ht���Z�-&0��E	���u*υw,���c-��Z�n�����H�uA&:�O-̒�a#�]hX��v��1_����Y>.�^C���DϪC':"�I� �dC�co;z:L���d"�P�������x�Z����yv �Q���D�߿�(��b��p���11^|Z������������=���ZN	[:�,�cƞ�X�i�5�%ô�*�&��܋��A��2EF{�M�=�z1�l}��Tt���S(8ѭ����&G�wr�X���ڏ����*�:_�=��hL�(-��`J�M��#���m��Z�M��N�h&c�#�:�ӿ�pϼ��j+bq� 9�_��bHr`��9sA�(���I��}(��H���Ęv�O3�0ةaϝnɟO٭G�,�Vw�)���n�q
���Ӈ��?U,;�_.栴>�?�i�"ec��H���K�,'Tv�����L�q�4е�R�i�-R��)���>H'���}�d2�#qe{AV�FV]����k<>�Gf�@���vwJ�d/��h1Ѥ�T�@����^�����E}ր���W���6ޥ�5��ʮڵ�{#��E���~-t��ʋ�x�#M�=��{g�I��ھ�m�b%4b��fg!��ׄ�u%�� $H���+p� A�I�	��7&bs�3z�M�UsE���f ��{��"�*�>1.d����\b7��r���^�w��� ��1�W4��J`���;ڑ7ʝ�Zt*H�]���p��H�:^o��V�q�F��Fu
a]����`#Ǔj��I7g����L�a#oM|�ʇ+t�G&Nm�+:o���m,Ȗ)�ٍz���SzBL�hgc��J���sD�Ђ:#��l �z�����������v��mg̭󡔑o ��L�5n���}O�JUk��R�9 ��
f	㯝4���0�0���� B��1yՁ,����Pi���1Ƥ�?�/�Xs	��*�/���9��q�A_**{j^)
`*����y�صk�R�D,��U8�X����#6�P��
�
2����-᠜HV���4�g$����̛yF��Z�|Y��1
�kp�#ղ:`��;�m?
7	y�H�L��~-=�x ���TCv�Ou�?���	vc�:hu�R7/�Ob��كv��<7�n��WS��/xm#?��8�,3����ψC�F󩖑�"!�5����݉$�3<s���~໌�%UdŨޑ�˱|�'x�u���n��~���6�Z��}�&�
�]�Y�>}Rp�1)p�N!D�9o@��!�5���;w��pL<�"�;��J��Y���87��\^Xe���h�(QF��v9�_كK�Pm��.V��	|+Z�)K��+��OQ�!�߶`⢤��IJ�c��!K`����0{�� k�������>w��\W�R�c?H�¸�����vtbߒ�T�Z�H�!ޮb3:�&r���}
=��a�+�|�T��<a�,�7!M�C/W�2���m�Ю�iv����m���^��g�c��-6���@����=u/�Ԋd���n�
��&Q�mr_9�����w[�a�)�f|������%�_�#�L�YQɌ�OW�N�3ԘC/��̆|
�<�å1��ٯjLea��
��߇Gπ$���B�t�㑁	�ނJ-Sbs��X+����O�x�r=f�2��D^�����9�{��FE���ȗ���n��O��՛�Y�	��n�^��ï(Q�f:w��!qLԤ�B)��'f@%�lKH9��u�aYYa��s���\9���a���d���W�6� �+��s�����4QBA�2J|1��:��v��Y�MU����i;���Ÿ�V���2VXQ$ӷ7��Y"UW��	�����P��% �(`��y(a�������c��l���TZ�H�r���E���;�$��1��jx>)=�l�vW�|��@�!1}?�I�t�D���p4�?w����ۘ8�_L(�m(��N�,�����>X�]����#.ĖG�0�0������O�O�M�q��(���(�J*�b^�
ǠY��/�emC��Q;jg�?ޜ?�����=��7	�by��O�� %��T(aI�� N�ߠs
S�릥�/,���W|27�v�1�(�_�͕�#(�tx��p�e�6d���u�C���)4�3.x�zS�.6R
�<�]�~�lm�����|��t�g�]�{"�|+�"�^��g'��#(jңH�B0v}EI_����^6�2�A_A܋����G)��/�0���`�a�%���V5T�6����L�����n�%5�xb��������b����qh�ݣ����C=Ŏ��|���-����ӑ%�؉5 ���w &Fٞk.�$�dٷ=Q�r@���F����ӏ��BA���ћ��@ؓ�����z\���Lfn�>>�ૻ��U<3@�$D^ؑ���PU��&M��T�	K"�DD᭰j�"�Aq+������#��H��UϏ�7H@H��mʯ]�<
0�x}1�8��S[�e7�*ݣ��	] ��j��C��j���%"9��M+a�����f.���';Ӡ��C�yO4�k�ato5���^����w{xbԦ5T+�Oޤw���օׄ��T�l��DlX�ܱ�9{��C�T�IgbAU�J�ԋ��_Z��d Xyr^[��b���
����8&uq�O�H��B̮���jdE<�h�Zn�=y�>�tX�N~��'؛`��&�:�IQ�Ӡrnn�)�ƝCn�em���*8	|�}�Y�6�/{��.HA�G?	��뻄�q�Dl&�h�y��~��;E���-_[�rYZ.�rD���qM����,�R�+�x�J�����E�惜D�C�,u�w�H��<;����u�1PRҀ�H���P���*�R���Ȳ���xe�ȉ>j�}0��G=�;�l���/�����Y "vk�r��B���~��c�(>��Ê��0.�z��!�����
�;�(-���:uhZ�����
s������>]s�����Ч�D��R�W-�� I?�
�Gci�r���@�t'�����$���մy�H�y�Uǉ2l���¾�{+�a�H����½1t�������P�.x!�F`N��봕:g��G�R����d��nZ�l�����#�Ͼ����n0�E�j�D��uͲ3, � d��V�s�Ç�H"�\Ŭ�5Y+�7c*�f�&�e�4�N����˩~D�o�W
oR͟��*+i�Y��b��^1���������@sg#��rA_