XlxV64EB    25d6     bd0Zj��Bj�s��#�?�nG(zU(�-?�d��DqX�.�Y5�tڭR,��2$���ը#5g{A�!d]��kVx�:Ɋx4��Knt����!�{n�mQ��r��ϖc�w��J'UP�3�&?�J���TR�Bld�_eѳP'9_KLq��H+�W�I�uO[3Iz�J�� x�Y����>期U�C�3^�^V�;��Z~u7����~G��^�\� ��H˧بu%�~�g2(~�/5tw��O�ڎ�4�}�ۙV[ߒ�X�]�˖�iM�X\�7���1���w3\�ev�����0��@���L]������B����^�P�0<�k-�h��$P���\f�R+6�,j�i�|P4u��x��%�~��d��SD����iQ���u�:�X��9��Hz�4���\��{, *���OL��D�휬I���\N�#:'�!������TqhQ;��D��,���M��h�J�Mֺ�p��c���~�B���i�q�Y���"e���]�Jl���~��5):����4'f�b����A�Hg�Q(�g���L�h������)A�R�l@7P�G�ĢN����w��]h._]�s�y�!:�I��!�p����nk!�S�<x�(�AJ���|����M�n���5,��U��epn�6RBG����=8w�v�D�TM7߀\���=�1�/�5�'�k��5!���RN��c��"%f�o����z��*�NdkOqA���^T��Ӷ�n`NЄ�90iA�_-ZZ�𸔰��R��G�����z̞3��;��yU`�i����]��K�|��_.����V���N�Z�oL�� j�vFd.ÿ~s�T$;����37���x.a����nU��X�Q����\r ����-Ra��DxK�qX_1�a����`�Ycɶ�`�͑�/��A�/ϊ�o��u�E_a�dBe���J+���T�S�O�a	%�)��x%�q"E�|�:�t�|��e������6yYh���0��ǌ�α�" ��D�J~�W=��C~JvF�3B�LF�ԥ8J��Px��+
����JJ���M?�M��?���dZ�#�eKlj� 9�'Z�L댦� �1:��:�� �B�z�2fsk����G�$� l�<�m�|?��u�(7����:;��������~����W����B$�"�	�+t;��ӗK�3\k� �tU�3�H!a���|Rg�#Z�#�|5��A����Fj1��"�Փ�8�2�|IhQ�� �x_��`�l[:GLI�L
��O�b�=�{B�R�׬j��s��<i�7�kk�EB9����枎���H��������T;b�q+
�/�j��e��U���x�g|Û|���D.W���$��z�p$U�s���Iz?~��V�=zh��c���?權u���[U�d��؟������cj�c�=N���H�(�7&���5�����i��~]XwEѷ��L>m��Π�����p�_���"K}.u[����ࡀ��ȃf׽�q4<#�t��.A�c�����(�P������!��� � ��F��ݸ��0��7i"���i.2+�m���_&�y���v�z��J���e�����NݛrO܍�af���+i�~!� v�Y��/��V��>�u:w�������y?���
�ᅱ��\�PD��o��Tm� |k�q�&2^J��'z��
������nvs��K���y�-"͐<C��3m�9{q��+�!S|�C�cdx�>��w��$��8��㼯پ�m��j�,�PW�����H��H�g�ܮ�Nq�b�0
5ZM�z�Gk%�g��8�׼�1<��'F�q".�&;�	�Z:�pm*�	����FSy7�L�]�4Q�:>B�1��B����YoHV�"
�aJZ��{�D��kql	fZ�B��1>�[=�^W���ښjCY��yk;�
e�9	��1/I{&~{* ���8
��=X���#�QedmQp��۷���8G����i-D�>L�K@�,��7�_��1N@��i�f�q�O��d�����Z3g�/��PZa̶ d��+l]�Z���
�Y�AƎ����jL,Y5���X����:.n��t����L�i?�"�����azm�f�F�{ZO��^K��꫉��oP+-��W�z�w�w佴vI��~���	�s�uD�UKU�.��.sI2`� ��.�jak��2!`�7�`u"�h��`�r�R��6Y�ĸF ����oda�~�c��]&��o�ik�Tyo�v#Y�=��E\��,���+����1�X��3�p��")@)h){�][��o��m��a���jFR�OH
mRU�?a�1� F^D�&�E0�b�Β��.��W&}_���o��(d�p,@}�7�\���]��I������^/���5�4�/��brߣ�3Q����+��m�Z2��ȭ�������/���$i��Zs�2§P��ů��k�I���7��є�z�tS�P̥�5#u�7 ��4T�$�����/Uz�/�-.Zih����#�^DjBD��na�g���= �}�˲H�㝮�"��Gc�`w�V����.P&��#6��B��F�Ϥ�xù�س���
�X����&jG��8t�+X���2(��0��s�,�����js爦L�(={��3DI}g��*�k�z=�E�Tl�4L8����,�r�k��v0�S�a^�0\c1���_���i�FCZɩ�ūC��b�PXt������D�R��@�F���ˇ��Ťq\��+�5�oi��ȋ5���V���ImWXo�Ґ����&��\q'�Ah|��m���v`��� Z6j���X��`%$b�п�KK�5#��%����,B�������7Ac�'�#�|�Pɪ�
H�Å�n�
R�����|�b����|����#ეx����Q��s����H�FDF[��ZG�����