XlxV64EB    1d20     9f0��WB��@:@|E��b���,b�:���J%#t������5M9�O�!��W��"����5�+��Ȇ�K4ػ��b�2����f��4f�33I�d/����+�3M�5�y@�syj
�>�Ŗ���HI��q�.��^�:��yG:%F�������Ҵ�M�����G�1��|��®{�Y��}�H�5�G���k��g��@(Ð��INr�EfY���Z����j���������HQ��u�,�w�fF9;�r�8��.�'9���;Q�uL�S��7�+�q�E��d�.�2�<71+�����{#i���J�o�ν�=����#ס{zݷ؜y�Y-��a���@�\�{�J��ҧƙ���&�Q65~FD�[�uΩ+�;��M��9s���&?/N"��KlX�ǻ�#F]��8�����f�f�{A�̼��Z�2���)�#D+m���A�6u-�(��~�+�H&[�+���%x��\5��A!S2�|ٍ�M�\C=+����E� Z� �~��,(}��v��Z�)�L�-N>��aJ��G��&4�^��)�"D���c�f�Ǟۨ	�%VEV�W&%x��*�u}���+B�t�~G0 7�*�E��z�)6-�Bƻ�n���R�B٠*�����2#�";�6n�S�=����K��Uh���յ�UԖ��\�y�� ��XUZ�H
��W�x��N&�uP��z��K�
�����+���ӫ��,�0��]2�.(��b��^��$�Cߍ���iJH��!\4Yk���:ƅ���A���LZ漐#�+�!�����U���\d����by�Ud�&�E��|�a�1�v`p�e���8 _u8�*�9ؔ�o�6C���cG�q�~����7������^Ā;��B�ڈYKu:�;%>b����4�g�}2���o;{�\V�飙��л!Y���D�{2�7��"!k6'b��҆�XX���E�>0zV<P�#������M7g2u�%.��yZ�d��(��z}X�@�	a����l���،�;�/���d��u�&��]�v��,���W��BY�Y���,�;����]u/��n(��2����x-��nb2w�� ����w���0�GF4�pۚ%	z�f�U��яC��Jw�T�Qb�N�i�� �6d/zj��9��~L�	gL�rF���Z�X� M���h��A�!�*�s��K�q��'�}|���;{��fY{��ޥ,�Lj:#����N�����s�Qp-�ۻr֨����Rk��y�֜��3m�m.�'��>)I�[Tn��'H��zo��Ν�ۼ譳�=�|7ŋ�
�V(8]T����t��6��؟;�.�Zi�hN^����Q��V���c^�d��M�jS��
V���	���]+ ������?ڷ<��c/Ѩ��!`��S�~(��J����o�c�"?�t"r�m~�*7��kH�r�Z4�-��?@�`݆� ��)��4C|W�`ч�����_�G> � �Qqli:����s��'��5�_�|�&x6Y��rY��;'�����{T	�5����!�ڹk��3���H0ܣ3Ln1k�J��{���De�6�ozi~;\Ϳ|�����q#e��/l����,T7�'��\C7������<��~�E�����-����q�}I��*E��]�X��f�,@p<
Bh ����~E�V�G;�g�:%��G�|*!x��0���h� ������ /�a�`J�+y3%,]my'%��C���"���D�q_�ק��)�CV���ۭ.�1�
C4��9DA*��(ߓd�������68_c+J�e}���@�>k�̺�ekUg2�U`XO����n￼#��&���>Ĉ߃��|�<��3��B��2,?$���D�}Z��ڀԒ��Y!�7�!9`q��j�U�W��63=�"u���Ֆ@�ȧ���ʃWߥ�IҘ��k:�t�����F2 \��qrJn�S<EC(��F�o$ ���eLd����د4���a�=8��[��b��!�Y��]x�˒v&��V��b2MN 1E�T$�C�5j�Q7�l����P�S&(��Z�d.0Ur.���t�`>�Ph�'��Z�0P��D����"�f���PH�a2b��V&���xv�|,G�И�֤����$�zv!��i}0L��o��:�Γ�:����Yn���Y�B�c�9;#ƫ��*Ew��s�GYצ� �ȨD�Z�H��l�0f�hvE':
�i���J�_5#!,�Pz���^�֗E�(��\��C��a���y� *<g����3�H��]���챑f����t��LŇ�e~a+�-������d)�T����T/��gI}��,�	Ȓ�T0N�z^�������<���ZyQr��8r�7�F�@�
��V��a��`f�������؀2���_ś��$/z�^6ܢ�(�v���6-�5/�ܒT���k{���(�!S��d