XlxV64EB    3b0f     f00�]2�d���b� !0�d6�^�QX�k�o���iEaD�O�Ǌ&aI֣�:^c���զ��׆�]}S�+�Nk�䀹=�2ϫ�I�!gFٙ�~��縝��[�(��ٻ���[3g��9�J���Se��lü�Њt�e�����X�b��^��C>57
֣��F�������5��V��J�2�16sq&��G�i�-\��O'G���Ta�<}���J�2��(��^ӹ�G�fل/�=�����P̏��)��i�^��:�	��Es��LO�o��Q�%��UZ8h��@ki��/�W�9hp G�P�T`�!m�o�'
!b�JX)��Y�1���d݇R&�H�4O�������A0{��"����
�ŧ]���r��/���pw��'A�£���C&�#jJ����<��q�xB� �?��c�:�L�x9��G2OC�=��Wz�Ouqgt�h7y�����fI"�o���5���T ��{\'9:��o5��9 2��%�(���y���M�'g%�҂ֈ����'O	-ͫa(��P��bn7��C^��bAh�Nb1w�=:ۖi]���⻥B��v%u,DF{]zN��7��/��nL���bTI�?�F-E@v�>\�ַ�J�ȱ�!�OL`'~6�^���v׺��$�ؘ�ԓm�췱|הmڢ�C|mg)�a
�Ģ�)�	/~���'���Xs+��v|��0��:�O=ۍ��kߢڌ��0���_�3|�1��7�N���3-a��Fo�E7^�'$^��ύ�h��@[�H|&B}�^*�՚on�7�i�|�Y��K�a��rG�6�����(�!�a>����� ������i�q���x�&ЬF��f���f�@�ٹ<"\cg�RO�Yb33��şTi1wM<К��έHoN�r�sX��]�x�����qٓp)D��W��-)�����<I_W҂ ��8 �[�_��8ndu��[�w@�ǵ4:VhN��:���B�����đdI�T���m���D��
����:�@�DZ��^iֲS���l2;|�R���؞�&�		|�HPrE�"Ӏ1�CZ��Hd��ƿ�~|s�6�A{rӀ"�D�� ����s�]j�-�Լ�Rϱ��;�����;gUO���ap1����ks�V��:�4ג����bUHv�	5�ew4h�7�p`��
�"�|	N9�K�ڦ��d�P&�0��F���,� j^!Hu��bkXE �׸�	WO��n��X����Ӿ���jY0�<�u�^=��#���F^�v����Ŧ�wao�0����Z=�\�(�3�V�F�fwm�q^����'dͤ�����Zㆩ}��͕s���5m�x~��*տ�l2D��G � �1Z]'Zcϔ����1��+�����۲�!'�#��wz�g~l�������EY�bq�ȥ0��p1��;�}v����ט�`,��
�M�쭉�𙯍�Z+V���E������v����:neӀ�:��2�,��}�����ꥪ_�4M�
�0��0��>�׾�JQX�f�o�V����|7p�>���w�}�ɨ��,�gU>_��Zp3 mZr�/�y����8 �'�굛�7!8����\=_��rr�"��f�lb�Ŝ&�ZT2ׅ�w�LϠ2��"��~��(�HL��ehּ �RH��,���Z��JO�u�i��%��Xǘ	a�2qp�<F��B��&�kda|�7���{� "_�o��!I+Lk�O������E&)j��+������Ӛ�'uǢ-Y�ź��I����^��5ud���J]8E\y*��/�f�x�4�����L�V�v�LRm���P"P�X�?���J~��w�%O'���&�_����Щ�EQXC���+��.wԫ�E�1�C~�o�I\�F!j��d��U���^km�it�4 �.@����Pq/�X)ƀ�����@dY<��kI������<ƀ?#H���� ������d�x��{��,8��Ƥ����̿�2,���9��%����xب4�:&r�jʄZ�2�rct��M�bWO/C�E
 �-%�aoI���4�I�˽��D�ểp�o�o�dV������D �-��yQ��� D ʴ������p�T�ͫ��dƊ�I
��ؽ�(m/W��Q�FH}IhH��!�9�=��f�ko�N�ğR�%���Z^$�}�gĻ����1:fU�]��9���j[�d��AtE���%QYFd�U ��I��8!��~�NM���B��6�r����_x�����,T�R.[�j�����V�}l��ܣA\a�,��L�j����a���˹.L�-~�D��E��Z�F�;A}xܞQ�BJ�
�ᶋLf�T���f����pa$F��s6��{c��'2�v�񬫉{{�c���=pp�DT9��9�q/�'���?a/%`k�f���Y�LW���5,껫���w���]�݋sc���|����t��@
_X�e+��K����$����4�f��P�'|ɷ<���ݵP�Br�h?��D}��T�I��c���h*^�����K�D����FH�cc_8�QW%����p��/����#m�+:�z��˫������ R�`�S�>�E?:�j<@���^F�'e�N`���z������;C�XJ)y�ړ$m���e:+������d������}B���t�Is�f�A�AU��H���V�I�����͓~�����H�/���防.��D��]��+2�D�*��H����I����{��K�w��A�C�B2E���)���bF�����vs��"�K��H�Ϩ�0E��&�����IT�'Q���b��"O���T|fg�ڨ�v�G��2l��D���u�-�'�B2#RF԰���ؚ�{����C����^5�F�DQ�Ks�Ö7ka����/��)�.���v��K�򙓨�.h�\dV�)CN6]����2�.ﵵ}���`�?�n����B���.�j�j�7���m�ʨ�A�N���b��W׳�Gx��E�AҊ��wQ�S{�$��;殲�AƇy�W�\��YS�1˛�$`�8�Ɲ�Ĕ����ў��Z&��U�N�z.�L4�9ҩ�L$��[���?�\�XY�cC�aIP(FG��v��#��nx����S���1d\p������Ӓ#�U�Z�w�-&�^��m�u��p��NmKdR��콑�Oܥ� �XE��e��/��"��E�g����[5O�!<&S�6+ѪJ�+H�RN�{�ǀ��Ó��gPʚ-i��#�CJ�ϒ�/�A��V4�ԑN?ph����Q��8R��S)��3-F��iK�:���rҎ��<@� �>'+�m��uU�T�����-����C���Q�Xd/��w?JF*.�����- )s�@�bv��g>s� ' Q^%���dj9�/���s��w����m
o.��\����7���8T�kX�|����N���xt4÷� ���(�gL)-��5�u1q��d�/��-�vn��ah�%�/Wrg��^�3�rhfP5o[�!.g�QL�u߉������ࡏ�A:�D~ F���Q����{��:�e��x�9���Y��)�0-v�b@�u�}}y�G�B�y{x*����f�׵¸���o���.�ϸ�\4 �Z6��m g6��(�ؖ��h�^B?A�V�Ҵ>����K�sNnԑ?�0C�9��ˍ�1NQ^@�T���$p'PAY|�ŢC�p-��,w�T�n,7�%�E�⹙����Y)d昋J�nPIߐ�Zxi�5
ņ�/&�*