XlxV64EB    fa00    2db0e��
���fYͅ�?9S	��XZd�It��V�7U�4?�y����=��y��M�D��ܔ_|M�{͹,��H#Z�{o�-�נ���(̇ͪ��g�T���ȔPЛs?�}-c݄o���y)AڢQ�Ǫf�#��:�̩���j�]��A�Yq��<v���K>\��N.ӂpo`SuP
٥j���8~{CV��ς	tPN���_H`x��-q���@��s���&�n�FH6�R�Z��蕡;}Y�m
F]:��H�ЭS��m-�8l ��/�s������Ѵd���#-�S`���$+����`Ӯ�(�r�\�>V�$<J�*9f�g#�.1�c��GM4�0G�u��p5����I,0d��{�D���!\�v�W�5"z��KI/>�g�& Hblaڶan+~Ʃc��Fb�����.Q&�ޣ���l	ȿ:�F��qD�&�r����� ��hS�����p�o!S0�Y�%N�՚�f1y��<�`Aô[�n��㿊S��|���<��h����{[I�6�Bج���*}���I3�h�y�Q^8}2��Ys?^\�|�ȳa�)�Z��Ʋ���$�v��;t�d���(�-]�4�EL����)�h��4�-ݺ	���Ejܜ6g�O.�d�h¦��빇�\�z��G�IX7G<<�Q�+z�;�l���B�4���j>>Ԥ�Nd�}�/�>��C��SM�;A�y�� �?��r�3�]����s|��)�F�s���Ѿ�⳻g������b,��������Q��BV�i�v�´�V��%�+�ڂ�-s��H��#-�w(�k�'�b5�����2I �j�
�IM>wu�DI�X j������|�����W���-X��eޏ�5��7�L2�Ӡ�qT��pMi��� W}X����0$qH��IEV)$� �6ޑ�QLW�	W��G۸���d�Pz���������(�C&B����}���|	SDpu�YK���e����8[��:n�=Cb9HZ�gd4�i�L݂F���f�V�����bc�?-���Y~FsL��x�IiW{��m��JZ������#W�������zO>ڶ4�W�iymT�'�!iש����U�_ٵD��V���	���*[��?7)>p�N�Qn7,�0x�DVʰ�W�8����XӮZF�HX�0�JAb�OS�`�I�d�=��r���%
��W\�E8��>q�T�s1��]f�� 
[�����c�G��� �Ԩ���ؕq\���r=X��ٸCQ0�.I��������QiW�A�!�q�, ������ð,"�_����A�����U-r��	2�sY��rU�ک?��Y���`ʃ*��Y��\� �r�fj����]�����a^��ON��\ P�^&��?c%h���ߦ��ʲY��w�F��p��N��I���m	,K��wu�jpnh4���|�, ��|�C�����j\��K;���<bG-� �YH#�^R�$��$��t��۫�G�@����V�{)v<�. �|R��XtE~C�]��eҦ1i�U :�y��������N�v%�����2e��	/S�G���S\��)VٿM�s�eĔ��O�~r��X �8Cwx\IF�`�YY�a�%P�3�ٞA1������t�-����S��B�BoZ�9������w4�2D���T4�:w�ͯ4�]�?�&�R��t�$�8��˃`�&�z���-�J�+�"VE�UI����O��H��蛐�j���)|s��D����e�����/09��q�Pǖ��
���m�q��^*�Q��"�ŃA@�q��,n�.Q�A(峫t�|��t�o\Bk�6�<�1��<.��������o���t���P+h�\	��i����*���ޮC�D�,hlO�"����0��Cy=Tc��0��ڂA�f��$Qe��x{[�"�\;�<��g>\�?����Z�V(\y��q�$�����w�Xr�z��"S!�L��n��΀�q� ���t���(�io5eRS�Y|�����eʧ�/n��t2���-s�������p��ɼ��4����9GÂ�M[P����w�E!Z11�����_��DV���2u���uWo�!��3���[�?��������"���#'p�j���Ő�኶w�y��c�1����U&}���E�:k�Yx�����'��W�����I娎�\�|J6�}�
C�C��CX�{>2FX,1V)�D9lb5b�+���ZI��o_^J��,�+X{-A=%FJ;�m���Ty1�q����(2�l&t8�������yEL�9��7�������L�JƲ���ݖ��<��~����"�Ę��ZFW�����5�J{�q�w�.���Yd�`�=1҆��:�$\NC}�炇饚�j�� ����G��4i��}��f��c4�@��>+��d*�,�)���W%15��\+r���{�_����$.{pW1�������o�[쨏K�z�{�Ih��T'%�zC��e�3�q���f\Y�R����n����t�6V�{��N0O��lH�"m��ŧ�%�ϧG��_�od���x�����"��f�|@ܹ�SSF��>�5��D� �������,��C�o4y?^'
m���τ� {�f�u?'��j����h�h|�P���W�8��Yi͈�P�kY�f���t
��_�r���l��9�&b�>�x�VyN��>���k�E���J2�=p��y�!ć�?� �`?��/:<��W!�:�<���4Jg���Z��=���%��}�ֲ��f��Q	a;-��"�8{n܊��'t���(V�4�*�؏�1����#�7فu��O|2�b�I����oǹKh»{ts�Ix��;�]�f##d�6��L,��W�c4�y�y��/eN5(G\��Ռ}�M�}.�S�)��uA�[���rr��Vo\Z��aUK�s��E7/���n�V]���h^�qf��l �M�-+&����g{Ԕ���'�@�	'�$?��Kb�g���#��_Hz��A�Wb��[���)ȍN�#	(>K?�?@WSf��L�wra#:&ݏ��M�Ɯ�$d��n!A��Jʌ��je<�������R�8=�)��3��i�z��	a�^�"�u7��nv�yy��:9<ܿ=�	�Z��%�HL~'W �q�F��x8�zT$z�<�r0�jc�&zu�-�\��c�r��#G��ĳ]�O.�:ιR�Sq(鲥�f��[\tB�]dHG� Οj9���To�(^DG��
մ4�7�u�x K2����z�+�������(ZϋŧWΚG�Q)�����պP�������q	���Cy~1��y`�y�-��G3��Aѡ{b(��4�������9B�2��X�/��z������y��D������"�+���3y���R�� ��aZ0H�~Ɩq��m�WjZ����Õ�/7�f����|P*9�S3�!y���U,�<���p�/(d^1��g� ,P=�jHM�	���+o����*M
�3��D����0�"|�d�hW{ZS`����>�i��.�.U�&����_(�PJD�90�@ߏ�m�|�/�v�׾��+]4�P+Dʋ���8��C* k�����
�c��E��}3#���@�v"�kF��Ug��۳��V�y�|A���oS�`��)�(g�ż�o:.�3��,����rcX>N�1�f5�=Ѵ���C��*�������*�H���M����C��� 1LvO�^_
 ����W*��
�i���f����R2<�~67�ЃV�#�� 8��x2�\On�nR�h�t�:�A��X���C0J��0&�����iiw1&�7�!�7��Y��_NN#���ZV����c�^�yg���P�^Ycu��2�5�>���1����pvnj>2���P�:�T�r��[9ٙN�I�2����ie�R.�.�+� �8dh�/wex�*g���j��9|s��#E�/2�ru��4i}�yK�%�9q��J/�v�0�:��M�韘- T@u��a	�״/w޹�-�;���y )6�b�*�l�qf����O��9��Z|Z�6�]HU�� ��'S6�igڃtx�[�{�D&M �ZW�`qC���h������� �+�眶ֱ�i��G!u�\nk+�V{V�'y����)�S�OY�ť0�+�.3��%�=\��?ڢ�
��j��"b�G��Oz�G��{����u���Es���A�S}��h��֐����Tp�/F�R
����������-m=�g0' ��z�꾮&qy 3��0E� ���ut�K/�8��5�.���i�R��c{��jN�H`F:a��c��=yu�$�K��>��೉�}fF�Y{�n�4��!	J�@����I��V�s^W�J�N
����<O�"*,%6B��������N���A�&4b�7#����I���$��ۨ����Є���I��3nD�"��NL���O���TlNs�@Ns�.�P��^Y����R��5�yZ�ؗ�$�{�s��}�Ԣ{��H�iOl8�5��Lx���5��_�ll��Qq};���sG�j̯�F�t2�^D<n+�8SR�U��(�
�c0뿉�{d��D�x��d{�٦�RԝK��xq8��Qն��|nK`>X���Gp�Ym�N��������S�.)�FI�`b�q��O4�/���s$���J���cB��g ��|�D:����f�6��#�	�۲WKi�����29�5���i�Ժ:���
-��6̠:�7������K��bf��s�k��v�s=����WR]R�'�|޵��c���f�#52��7�91No+��& 2�E�1��E��?�sRY#�7+@2�:Dϐ���}��U��,��
ь~6�҉ǀ�RМ��cݠv{	�(��g�n_@:��K���o�V�F���䂡�ZfR��T�G�����[�����XF�}P�/���t�k�,RA�FomP�c��{:a�6�SW�+��y��-�8@���e�~D��c�lI�K��Y�S}�8/]�WI.�G�wZW&�Օ��yƩ��>O�t������K{t�<���}�r��tV�0}�����Hz�(S(^���:�6F�7xz� �T� ���Yc _	�g@�W
ݡ_��*��j���\,$6��������H��S��.�h��yRv��>�CO��������iS[؋C�|�*����ѻ��Wʲ�G�(o�d~
;�'A�(T>���p<�i�Xߴ�͵�b�/W��|O&
�ó����'�2B;p�HS�C�Y����q��o|�&��m��
:�J��"�J��`
?��@*�Җ�*!����p-�%0���
zO.����8hT�y'�W�2��oK�t�TGN$�#�_��$l t� D8u��$��~C��Z��
{���mj�q�z����e�jZ>�N]aA�WDjO��;ُ}��w�������^����̙b��m �L���Z]�-(�S����1R��T�0|1\;W��7���))�m"�Q�2���7�ϐ��i�z�'vgER���X���5��z�8���'�3T���N�C�����T(��å�Ӆ4|�����FE�W�ϋ �Bŏ�������ڢ���`4�+2
���3�O��l��=)�gI��v�07G��$�=��J��R2�{�n�5�R� '}B�jZF�P:�|�"�`�|~�2�������
��UQEaU�:z�"qq�������ϋ�*�{�M��Q6=��I"�����0b��_�l<������2���P�;����t��S�T���TT
���h�s,W�&�6��hu�Y��ڴZ��D��S�ql0]���ڝ��jb�d���e��C����5����b�$�E����M�_M��`��g<��	��Ni�v���lχW��®>���ˁX�êE����������J�;�8{�є��<��m�ɲ�#l�g!��v�P�p"E��E�4p{����>���E�t��BO`�+�b�"H�-�KF�1Q��������� �R��{�)1��<�,$��ʴ�uF��u֣57�(j��p����B&m�G�d��cv�W�%�>l�{�g�s`!�|�N��:v+�#=�ݳ�~������c�H�"f�	T��C� �ʀp�i@L�@��u��]Y�K��J9E��|�Z�:`��'i*��y������vޅ�d�uA��&ޡ������$�`v�A���9��J[{����L�s��O"���i��X�4+<�v�F���~��7��&���nAc�%î�+�n����i:��|�2��U�� Kv��L|C�OK<�,�z
�>ȲB�BAED N�C^_������X�"5ܔ6	:����r�v��Vu �x�]�[l�@��W���qQ`����n�^$'������V�d���&��I�f�>��� �3�w,��l��aN�ڐ�����|�=n�ĉ!F\1�t�.�[�J3��?�y1Χ�2�X�W2&3�=�Z�������!.ZE�����?�p��+g"�M�೬�|�"�?Le�"��c�:��_�G��V�v�^C�� ��t�E�rl#(�.���1O��0�o)?���T�G�f50�n@U$o��a]�b�W?%�?��G�k�њ���� I��3�v�/>�9ras��>k2DB��;���ݽ+����>����R^�UNħ�'��~������KA���-=�]�\��?|�!8������j���P�>�$uW&����i�#�ys^���fǦ�o1�$���ez3� F`�@��]� �=P;��I���T/;�����͗On��o[>@gש����^_������i�P��~�,#������n{؝2��OG�p9����x���P�+��{߄�la���q�IP%|��8S�@HF����_Ѫ����oXS����ʩ�D�xPuۭ�j� dP�}GD�;�M��c�GNҁn4uY�b���xHQ�5�랑r �M�y.�%c��U|GfX��"��%Ia�M�o�Ӯ^,k�f������F��w~.^:�*e~U � Z��x?��M67Wgk�C� ����,��B��	*gI-"{2C�c�����6��KJ{�_xK�X�Ǧ�������5(&��0���.�4��	�|$����̒��,rJ��W�´M���z��䔓g��OA�2o^�Q'`g<��dh�K�T	�R�n��';9h�l%�HG�icëur��A���Cb�3�4�z.��R�y6&7����l��J�iim��ѻ��y��.��-�U�-��79A�]�U���J�mӄ�_�t&�t��|��u���&��ʋ�!b=�%�/�{$�bzE���;y������h�C7L�}����O�p�� �SȊ�D���?aG��U�^��	V���VY(\�6�W���鼜����A6����+:��>�<�ӷd���B/�w�/�pg�����NĄ�L��D
	�zN>�4�u���*�����nD�d
�@ϲ��H$� k}z��+�C���$�����<��a���˿_�����D+�\��&5�f�Q��|�b�ژ���HLc���O>H��6�E3S�*�H��4?�^D$�B"@���V�}���$�e���2�*a�{�� �s�������J��m�,���L�&OR@�@��/��fӏ�UX"����%Φ�bl%I�fyG������
@�J}��Z������߻*�S��L�����;eE����]���x��q)��9\X�E�0*#�G7�U�K��_�����*�����!�����֙Qr�^�;"wǷ�zD�VJG��6c�/����X��l{��o�?�%!~J���}ޞ�����=!�u~�K��`)��\:d��>�I(� ��W#���	�e�߸꼭��l�j��A\ק�0�@�{���W�_wl�	y�]����dL�`���%9���u���H�ǎ<�+��nb���y�6Q�a#'���r�;��i�%����(}�Blw��WSq� �M�Y����
��c��mh�z�p�b���N���<+��>	k�����(w�x�6�����m�}�] �c�	H[��u�vb�[��������S{�:9�o����5~�Z�WZ�Mz���gA3�%�F:�%�^���@p�/͑�B�P>���Cj������;���
?I���x��В-g�B�Gf�,.ߟ�c�S�nؕ�)��d�1k���g�<:��Y\�c�[3��fV��/߃c�����ZE(�	=��7��Mh-7����&Y�7b=u����ơ�H���v�m�k��[X*�6wh�!��)$Ԋ���k�U5,��w��u\ d�,�����K���Nm.M�H�e���L�.�Z�?A��/�ȷ�����2M�f��XjY������n��qێ���I��>�f.�q�L��Ǝ}�9��v�*�YT[tܧ���j��3ws#+7��U� C��
�+P ����Q���j@K�B�o�/�˂�@��N�.n��S���;�/�`,�cg>�G�P��T�b,:���,�Hm�T�>�'=[8?R("��.{���b�'���* O��'WyȖ/�H|W�В��rϭ�Mw�J�{�3���3�:o�q&�K7F�Ω;~1^�3,c�ق<\�JJ�a���� \gKvr�AE���R��U��dK�`|�ԛ�6P<hI�q׼��cK�����Y��e"�G�|+S\i�x�B<_9��*K�wb�g}Ԥ��m����ǔ�1����u��n���K�,�_���Ǭma��8�gy�?x�|��[�7I����wQѝnއ�5�Y�<��0��jD��ƢHRʴ��}(q_��c=(3�I��)_]�+f�hft����C�=�J�{���,{��N�gI��"Aޢ;���oY��ܲ~�i��������Fl2}ʝ�~/�����T�4�{��n<4ъ�� ��F~N�~�����PW���I���T���;Vlp��=Q�z�c�����%��Da�����0x{[r�ڡ����o�4ooC�zh[޹����z���*DS�It�K�U�M%<e?��5SiL�%�,�d����*orVRZ̠�Av���U����� ��Yi�F���|� �����i(�&���������j9�(��mz)HG�z<�.��	��UTo����`�����n����q��z�%F~3���]�B;a�;f���]�3@2����y��fE� ��|ҋ��ze[y�O`@��a?�v'��e�ౕN�M����F�030q���c�?	�j.��B����J�^k�1���TG%����(%OL�m(��R��V?
�S��<ĳi�p��~ ?�8��/<i)Mt����g.�4Q9^G_��AG��qw�G�.�|v���U#і�%=�)+��Y�A�< ��`�o�[�[)W�D��&R[�8���$��7@�����>�I"�'|����ғ���x��y�b����I�{o���~%�����lS��@&0{v���h�ۡʐ} �w��n�b}� �Q^�8�)�L�Qx��|�ck��X^�q/먻{�i�͇}���¦��g䝍�@�,�0�8N����Q� ��a@��d#1G�k������=��BR)�T�?x���.~k$f�;[�B/w� xۆP��ℴq�q�(&�����!qj�7E�.��Ͱ/h3��E|K���K:�X�Sy;R�9����`U��6$���r"=����U�>�Δ�'��|Hy_�Pjd��dS>&��=e؏]^e�Mze�M�i������[ER��[B�>�J�@Ð�t�Fq�
$���>h�5��*I�q����3&�h������rp���ƀUs�4H9+�jSz���ytL��>�b�a�<�jߋ�E_���j���wm������xI�K���L��gY�Ry��GX���4������[Z���9�����M�yfYK`n��c����7򷔢���|N"��9��xn��62�	��i�%lSr�����I�z�&��~�O����c�F�6���U=/Y�i��D�\Ye�'h��LU�Heo6�C�^T:�8�'���
"��1��O��1���-8��C��"Ո��ȳ2��Ɯ�k�yzk
A�S�{��߭V'-s��E��,���o1����8r�ӖC�|�^�˻�l���"���g��6���}
���X���Cu���n@��	z?7rǑ��?�(�ux�lb�j���TA�e�)�O�VY�������$=4o��-)ϙ�w%Ao9	��2}������{���y[0���cq
q��eﳾ~�O��(:�H�*M[�;��{�����/�|�������,`����D'�� �Y4a��*;��_�(�D��;�.DM�����^��� JRA��,+2�8�u�b�k��171�咊�Mf�>���<la�ZƆ-ؗ!YB�a����#����踒�s2��3��8�-��U��k+�{6{L�U��	F�O�����-}7@;�@Ym|����M��3iZ*�W3	 a�s"1�ފ*�4�5b�C�4��1�)_4��%)�� BNd��%yG�'�w�lN�\������/�p���w2�
�c-��3P�����:�І�V����`��Y��T��`_����,��.V5����.xfX�����"��C]V�J":��C&�D��x��7�Ux(�~��e�)^�p���Ջ"<J�N��O)��Q`9����o(�3� g,i�����cw^��\qpCJi�<��+�el�Y)���fL��P�lżJ�����첑FF#�4tڡ��~���4���ᒡ�D ���e	p�<[ۭ�q�״}��my�[֧� ���?��;v�DN��!�WX�i���r$r*uykiV�� ��U�x�!��k�V��@bdU]^.W��DQ����R�r�n�����V�·�[�R�D�_��//�z{�A�tf��p�nģC"x�;����4��R�vo�>S����m&�P�OC�&zǲPsW����;�g��{�?c;1�-,�vM��� @t<U�	=\��X�1��j�\/O�Ǒ�@%FY��zW��>��ҫ�M�z�"�? `ʺ�󴊊M, {18<5w�N}z(N��~ٶ�d�&�g�f���Ш�Tg�l ��ck��bh��6l�*9����Ut�p'���V��WX���$�lEz���/�6w�Ԓ\ǜʬn�}�W���y��{�g�vy֙�@� k��� �y��z��s���m1(�� X1�}9���M�FP�U�ٍ�_�Vo��U����2s�'��)���,�4i�#�p��3��Q�=���<�#s�Eo�u���� 8�*�Z��~���+�sv1����϶�oPGG���^����	�=�� �����/�*�XlxV64EB    31e5     930�UbW��%���eq;���O7�g���<��=�8��3	�{ۢ���Wʡ���_�J�|�3��W��0su(�A:\��CIR�ދ-�bM�d/�:Rj�2@�F4�2.�Y���h8W���w4��R�d8���I�������S���5�����e���e��`���j��r[Do�]��Hs��ŝL����)����o�PD	�ςW@5"��LeaK��o ��PIW��}����#��&����j����l������x�:ikb��.������n����ò@���\ǩ���� ��I��ٷ�y�O�{#���ة��8���!BH��ŀ�9����uܑ�i�f�|�,ו>9J���ݙ����#�a}�lP��i�
F3���TD������3(f֟wE��Q��v��Im>���LT
,���p�lGh ���B[��\I�朗��lF��c�ټ �g�b�B�w���1\�}c����6&	'ESza"���e�c�񢊖,��(��tæo(�N2���L�,�rro�5[}6o�k�����KD��B����m���p`҂���<ufz��k�r�$Z�;�t$Y���j!��T]���뼤��T�DD�]�),�V�n�J�I��
o�l�����D�.�T�S�|�����)����V�@�9�����r \c=��[d��E;'x:��?|��w:+��א1hK�<�n�Qe�7ql��m֗nfN%V�Q�����Q���yIz0Ug��UT�y�큺�4>��כ� �7X>��&����
��#X�>(w�괌�[6*����O�Z\�Dd���3�w��KD�Fm,�ܨ�&��2��45:|�m��8��:}�)�� e��2�|˫��܀v��F�z�z8�AK���i���=�"��������zM
-��nT�!���Y��+���џ���D������P��2�-E|�L�rG�W�->Ax�	N�x@�t%��ַ|y�6T�Cn���8����g�ʤ�*Ls'��^���w�ND}f*!�G���)q*e��[��N� }q�G-M0!�fzG���L���`�`#$���B�n�F�P�CK6�_ <Z�J��ҋD�#<�G��w_T��i[�>���*i�^.�~J���}�a�%)V�&�� �8u�e�@�#;���9dO�7>�/Q�d�j�� �>_�PP�!l/c��ɇ*�锰�J!����C�}��R�a�W�ܔ������`b��P�Ǡ�
�@�ћ��2��H)�Gs�{��.r�9j�[�bi�>O���J�6m8���M�>����'�)Svw�Y����a��(�ȝ��e�ʂ�j5"*�D?@���ϰ!c�Xkz���i�vŠ��t��G�YH���֝ 2����;�v���f��>��6t
��y�~��xd�B ��t�%-��	 C���&Ч��3�㷬�"l�Bj��|1���
�qb�t-��o���;!���,1�`�j�%^�h
�$���̬�	`oR)�B����bd"^�T�I,�PSc�$v�Ne�>�`?d�L�|ݠ�վL���?>Ji:b�~r%a���~a�y��3���z�-���4����Ay]]�D!|�����c�����H�Xʬ�+�]B��EǊ�qy~���ءվ�Q��O�FࢮYG��AaN��:�`Ơhr�}�X=�N�R�[FOB2@���Ƅщq�=a�WmG���ʑ,�����FȪo�����yh/��#��i��h�s���$��!��yh
�]G��q��"��W/Sm[C��B�Hnu�P���8�R�\�2hZ�e��8���-��Ћ`Uj��*!�����&~�]k��)�.O5�G��й��������	;I+1�G��H��s(����+~�B6������?M��Qh��]BOј�G_�aQݤH��bv\�S;b�(U��<�-��!Dm籑�;��0����0�2$\��:A��y�pC�@�α'�	�;�9k+��p։��o��?�֮���)�1�mʷG�����;l���������A�A����-�ņ�"7A���\�Y��'�J�
��}S����ҩ�۪��6t�I��p�������hPXd!']Xu �����~�./s�M��6�a4�#�tei�H�����j[��dW�&����֮�ߺ��1>cq23ui:.�����B�k´5xK�8E��x��WG��ª���퇉���r'�$ ����ax糠��������d�cI���q��a�rd��>��6;���4�0&