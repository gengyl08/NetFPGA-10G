XlxV64EB    15be     810�^y�S�/8)N��C�x���d��3p悍yp<��dUńJ&/����y�:����!=����|�7jp��c����wf�C+Zc��y�=��mc�4��S��2�uW���`{m����'M���Ud{�R��t��\��8��P1 T��/�po�a��M�sQw��7�CWmߜ�Q	�>�M��C�����,^�j g����i�g�LH u���z����hB��G���Jވ/�����J��%9�u���d!_�o���0I����^d���:��d[	0�5 �܂�ޝ�-�}�|S����Z= ����5���;�Kҭa��<k���=hH�e8��
�����J�-�#���n�a�Z��)����^�B�cg��g�2�������Z��g���LS�iq'����|=:G<c,�|����G.���R�JU�S���6�M��j�_jy(����y'�H�D�y��${]i��
���PR�;�:ř#�sw�AS���@m7^��=ǂx�t�$�א�97Y�!�f��
Jϐ�l��ƅ%H<3D�޳��;̮h�]�T_H�~YH\����b�-�<E�'�^sS�PF�i���Kg�Aq�����͋MH�Yx�k�������Go?V�~���7J��E#�g��0�[TN�dld�&��l�s�,�}�%D$Kx1Va� �qօ�<��9,Ó�
�O%��1�8�\���GxN��YEv�8O'��'f;2�$�d>H
$�I���◙R��K���B�|�2mBwJк��Jz>n��"��AĈ-`��Z)&^�z�j�C��S��:e��9���{	&D5$yܢ�ޯ�d�AënR��.�1�����* �Tw(:y�Y�FLs,>��k���L����a������;|8�%bL�����`9hWa�&�������)9�BR�
�d�A�Вң��N���oc���9��QcI�d~�Z�ˋ����\xF-�N5w�M����?��W���>�=�ҟJ*�V���c��F����(�I�ګ9~�Gv�崤�KfN#1M��4AD��
����qHȿ��y7�����3����(�,�~E�9C,nM��/t��G|�w��5��5F,����Ϭ8�É�\���"w:g~?��6�	��&D4:�U7�\�'�!E-�>w����ǟ�:E��������lt�S�bie,�@�tވ������K�A�f���K�+:����ӕv�v��U}T@����CF�����p�ƐH��p6���1�v��|G���m|��~�7�L%��	�����l��5���w󙺻M�R�vB�"}*̭-�j�y�B����~�߼\����4������T�2P��1O)�#�d��Yf�������+t282�\X-˄�t)��D�%�m�@���	�N6Ix���U��l?X,ZM���Qa:�ԏ��p�	��!������Aw���A*R�+mY�n-�?nM�Z�7f-�3���u�.�P����o�Q����3���x��j�ICöWL���%y�+5��H�����©�2	��(mp	K���lЏ�C��ɧ�6/��nܭz�-�&�^[�����P��,�����V�� �ټ*��q��3�i~��
���}w�ײ��;&��r�AM�npO��@tjso�ڏ�DO�U�H�ˎ3 ���e��P��oxx.�P�{���d�?~Ci%I����
�L�$a�3ѫ͢;f��#_��[���r��h�5
{��>�����)�Iݢi�U����͡3�Q�Z��Rp@&��>��v��}��h���"o�M\шXN��L�����H��z�7E��T�4����z3R�O~�ۤ&f����iTu<kR��١���+=��Ӊ+g�sEv�a�y����"�>�����$��W3����ixސ�;$<���_�M,
���?'�!��<ϝ�cը��b�����A����`��$S�������� Lq�"���9�9��s�*}�����]�V=�{��t��K����_��/�2�T