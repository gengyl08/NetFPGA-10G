XlxV64EB    1569     850�r��q��>�E�bW��cp%!r�y�c����`��k���O�K�k��^v4��Jf�
^v�\������'�]Rv�XZ$�7k�|�2<�����Ӓ�b\f����e�������th�w�C�՟*��a�@�iy�=�ҙ��ނ���V�y"�\M�ϟ��[)wCܛ=�?�?��`����G�?XH� �?;r�񓑝ѝ�x��v�n�)^���*���E��2gB
$� Z��բl|G5���7)��4�=#h��x����g�j��)ݲ)G��n��p�4�]x�� �:�u�}V��_m��i�m���T�ٌ�N�U�t�u���`)7{����!oΥ˟y~ܕ��a��=�xk�ۭ�]��J褯Vz���I�ꆼh�Нv�UI�M2����b>I/���9+>o�~�Li+
f�}`�����|vEc�dZUsҳ<>���]�e�$���=�c<�K��#�h_�[����A��)[�ȗ�r��3��A7���^����:x�����!�#���0����ve��<'��h��R��h�p���(���>�	\򆠷x���U�.1�ަ�6��1p��w�>��k�^&u5	O_E��zJ�7����l[v�`M�+0�HرYO?�zأ�]vV%���i�ncЕӭ�
4g����[�L���/��+װ��%*Bv�F K�~UIc
e�D�Q��������9jY$Y��<�)MH"�����GECmZ�yX�.Sկ���F�@PW@��[���H��M�4د[�ps�ʎ^ٙM_m����7�M'��9�١��H���c��F�	j�� +��������P,���5�GO�A/��v)��!�-����	���,�������: /�1��(I�l�11�q���������yH��Vw��.
ſ�����ϼ],24uqX���},�p)c�'�Qm.�1�&-����S0%��'S]�G���%ͨ ;M�(7��w��&�a��^a��Ҡũ���A�o�����������p�H��-��ʡFhÝ7A
����w��$��l��=Qv͏�#��@�c���U29Iʣ�����܄��;л��.$'����(����6@�l�f�,���%���X��R��	�k��˫="�Z�Н��Oѽ�@z`q�Àd#��B��Q��9���k�B+ �S^]���ަ-�[�z��ԗ�/\���6խ]6�E��ϰ=���c9�@M[C�����'c2�ې��J����ạr�'�f��$ܟ�[T��:I-��u+��W1��3���q3���̹���{Y�3��]�����Z�,�'(kG�s2,���
\����%���cE'Y��g֨��:�(n����ԅ��*�F`�t�=�'�;���B�↰�
2�e~W�'K��嶺������$���mޔ��+ˣ^~��5$p�e�w����;�u[XN�9�ҙ4\B�/6��fcY�ښ4�mXDU�7�+����W
u����#��/�Y/I���`�<�1N@-��^�W#A��F$��"U%�9�A�>�H
��\�b�f���ݍ�xn�ѐ����j���,�`�q�(@�e��4�s9G��g>K�_��g��e��4UM���OmN1�)ː���a(���Nkd!~y8lu�	M���M�Fb��ɀSr�5]�ت\PgV��t���ʙV�-Q^�Z5�:��p<t�9�ǯ�r�Y�x���(J��J�Y�����X�ɣo^�'���� kϝԱ�4�P�����se���7����Z$&��G���t!v�j��|"z�)+}/��R�3�S���pk�(,����C�ɮ̗��K,p�ɀRn�f��?��W8M�œP������{�m����I�Nf�j;�ZB�x����}NN�u5��&�w��e"m��`�8���l��L��H/<�;�r�1L�Wp_�>� >Z+	K�{�F0��1�!� ����`*�AZ��]�b2�}�!g�(fI6�1��k�A�%��}v^�V��*�HH-���4�VlLq��$݋%�^w`���|Y}��.䖅Fz((�%p�qR���AיTc[Y~6��