XlxV64EB    589f    1210�<4�bj�瘮� [����С�S��7I�6��Ɵ���4q��pw?o\��0 �pMA�S�au͸��_�`�+8��
(�/�>��"t�.$��ժ�L��^�u����P�ܜ�<�W�n%~��E����n��Da���Ub�*·����b`+�!v~F�Z���5My���������W%�����`_t�$ȞW����ۺ�I���ʐ�=��§�މ��_~�Y�U��˯�`�v�ӓ��r��E}i�!�Yh�*������w�u���(L��`�Q��|���'O�U��q��bfl/��V,�X���-��Y��+m��e��^�x�LCrp�A��W<�R�p��᭏�5���%3Җ<z{,K̴<"x���w��f�N����EG��[������͐JȐ��43x��6�^��ٟ�<\�8C��é�=j4�rXGu�Yd��;�2�9{JmS�۲ښ�YS��~���� ���Ai%��#th��؊�_�hO��mx�j�\qw逗 �H8�;˕�r{���������S.��^}O7h�_�9�zh{��.�8�6�P!�CCF٠�wS�>e	�SKX<���p��w��Ar4��n�TĊ�B��<jQ4����$�n�;[l���$���M4�r ll+rУ��'�ޠ-�č�gqMq`��6o,+ˁ�ӓ�-am�.�dأ���!u���l�7�|�>#����<c��*��c�ݛ(��XI��q�3rF �QwF�Xh�z���5���=�y�>��S
R����x ��]�s��(�~2�˫�k�=�MQ���3"�G�3rq�=�ڇ�z�l����B(�H�:����P+M���@���k�фД,�MGP���-���&U2�N;�^� �O�Y�b_&�ג��q�G�̤��O��έ	xʯ����Cʌ
=�g�.��)�?eM��uh�����C���"���%֎rʤq�����$�I(}�����x"���&[y�1#���{����S��GF(�KlJ�`���D��ť�b��5ػ�csݢ\h��>��xt���`� �F���v��˩������Tgu���%��3%%�dڋ2n��NuU������Z�v��%7 d��E�P�µ�J�Ͽ�X�`g��Ow�����pV���n�FW[|;^��QE�Q��� J��ȵ�I-�f_H���X̓r�fh��H������D�![;@=���?G��xkoI̤7=/�!'ZJ0�d9�;$#��j�+������p����Vq��c����y~㈜� �y�!99c3jނ���-"EJ͂T-@Aszz�`�;nL�w���&�s�E>�!vcl*�SmD(`��?�:7[���\q��C?&�ɲ����#�\�ZI�-���j�ㄜ�T�uyN[��D1O ˒�ZE����H��|�~"�it�2��>:���dl%���
���L�>+�w���}�ԺP���̣�mǾ>g+��l��Q��Σ^ý}a7�	�Z@�rtϐ�euνƾZ(j���� ��60T�9nYt��̕�W~�O��{���]3�Ǎ���eqv�V�?)��I3�?͌-�S�������:С��'t4�:³�f����f"��@�r��e� ��e�a�'�����U��I������Jm����"�BJ�0�%//��p�(M�BM�tm:/�Tn[�Ո�;l0���c? ty*��'����r=�a�p��
NQm]h�+��Y�V�ѻ�������C�G�+"Ҙ}�dX�!n��m��M��Tfڠ��a\�Q0�۽v�^��s� �ՃKy������R�D2QZ����ի��h�E6?-ۆ�c���a���1�
 =���,]j�p�1�&��:Y���/�EtE����H�F��ۡ@�9	$�&��[C�D��)�Z�x����7��� s�jFoF@�k����Ç��B��aʀsw��I������GC���_Zd��M��m�8(�lGkVȰ�/�!��˯ �)����� ΡMw�'��$�$�uy'K{]�����JM�&��=�M��O�o&�]jW}����@�G���9nDa�?t��a��&�-{��R����f��Z�*?p�3� �@>���f&�H^)�q�j?���<>_*uh���J7t���J�>���x��5�>K`��3�����4ľ
f��*;KI����N򯒺�I2�^}"<h�n3�7�Y�؍�2�T����RvM�!N*pB��b����]_�)D˕C�	�k1�:���+Ql�&F��C���X'�n�
4i8T���+�"�̭R }�d�c�N��\�H�/aU��W|����F���jZ�iV�L����`���^�7��H����qX�>����v+���_�i�f�\�j���p��G)K��k\�Z���r��L��)-W���	��Ԇ0Ι˺e�h���!�"�����.\]ӯm�ON�[��p�˚��i��BBV��#���\��&�/����m�Ɨ��ecv��Ԧ���?��r�fg��8�^_|y�4�@����ع��q`h[����$�9�(��*��F8�7��J�ʞ!�>nm�z��� �iI���qWѾ�-0�7OXAkx�Aަ�4��/Z;�ؑ�N�L�va)i�Ÿ:D�	�!+<�:��2�c�ֵmvM"������y׻����we�-96�E8�}(w7G��c��T(+���b���	O�"�ّ����fC&��o��K왗i��K)�ԥ%���5d�����t�USi��Z�c:�&�A*���%8�g�#t�D�%��0�^ea/=*
w��f���C1�tkRİ��{��*<nR��:����N�p�lbV+nj���ع��x�Q�� �V߈68�Dq_
��,�w�aB�uk�ζ�Ǫ?���e����:�1���F�U�`qp������6�[���5aO�ш�_/^�#��|/�`
O��_�h��zg���/�.�������V��f����=�0Lb��Ɏ	���z���e�$�����s��������6�"��
�F��/'��4�����W�lNh����k��������e�ZRVhن	= ��ѻĺ�1M��P����>�OiA+YQ_x�-[EU��"m��	������7WM�Q.D��'^^�W*nJ�G��#��Nui&E��I��茞� �W�[�"i[�����	m�_({L2ౌ�ET�,&��qn�a���eN�:/��'�9���DP��Q���Aj�5����X�P��+��s�<��;��fa��j��d�؞�8K�s?�:Q��[M�w\���~ۤ�!�PJ���YT,g�D���4i1V�Ħ��{I��E���Qdh��]H�S���"`�A����3�p`�,�cs~�.wo�@iCV�����bZd���;��Z�ޘ��*f�Z�x���:U�i2�L��}��[���n�~���!�r�kC����(�x^�h��k�NCJѨ�wR�q'h��9(5?��%��+'ip�e3B�~����g�,�f0�	�L�#qs@���\>xc��V�2����xR�#�u$�����߱&F:�|�%��N/�mթw�ʘW �!���o\skK$l@ŋ�Wq9�/lL���v���]�K�����B�L�3@�?��uֻ�m_���Z�������a�F=-�xN��P�^�����a�J؄������.iO��8]X�AE �m`j@zZ�"����s98L�?�J�p�w�Jfr����ŪÐOy�f(M��Ey�=�Z����;}= {V������W�&Q��P�!j��a�p���R����k�AQ��]�t�JU��7�޿$���@����P[frDz'RH׎��f�����e<��]t<x��i+1PNtw�N�{N�A��7��%�!�1��T��6�:��S�N�[7s�&��-F����jպx�nx�dO矪�d��g�TF�~Ԯ�[�,�1�9G�/Y�����cG>2��X���`�4�CX�'�Ąw�kM���wK��.H�>��Ƞ���7^=I;3��d�
�W탛��z����z���gB�ʯ�?YU�~�����=f�e��M����C4����~�=a#:sh\�&����rC�l|!8]9<Pe���T�rb� G�b�1���C4t��M�3�K$y��t��>>��C;76| N[Wc P�N�</�V���[�b�!�ռ���l�*;)��/��}�P�$�O
L�%3����q�:& �_���!g9Q�6	�e��sT1&���f"e{@t�BΎs����n~Hc��G(�Ų��"|�GB#����R.t#��̝�5VK�&:���	uP~D�zS���ow�O0��jDi���L�oV�\[��	��4�]��	Z���g���Qs�lB� V
2ܢ--��W�0Q��l^R5�?7�F���_�.���ek�?�`.[e�����&��D���qCx�(������##e�2h��:6���&XN_B^��a�&dXj�k�