XlxV64EB    7c32    16f0F�,����k���KD���ګ����'��/-��h���S�M{p�L�����\rQ����Y
�AQ��u=h#DL�xs�)�W�8H꿭2��U�Wl�V��1/O�p�]T��Q�^��2��HG�QGWj�Q�{q�Μ����Z���+0�N����;+���+�q�S+����1Pcӎ��
?�1��GUu���޶o�|��ݜ��-��/��u����f�
�E�
�wY�b�~e�Q���H�hJc���T���G�+�9�8����7�&�x�
e\o��!���|E�+���
N���_�f>d$;�A�-؋�MM�FCT�
0a�ldc`�P�l��7Ú��h�����n;t�c���kj�bk%��Gw�x��C&wR���l���8e/id@�0�U���Wl[�=f)v{�.��88�C�U����Ǵ�b
��I'�RN	�wuH�Ӱ�_i�v.��ԫ�������_�����E/���@/ۨє*lO �?��a:}\C�����P� 	`�7��.S�"j��E��j\�:v�+�?v�Ĺ����l�0�����x�S��68����ע��*v���\��Z�lB��U����M�AJ��"d�ᷱtI.��鵢IN~��M �	��ژ�T�p�4���c�X�.=��U�Ẓ����k�F��
�i!@����Z�����G8���D�����TUC,��t���jƅu&�{�E��q�+�������7p����X2�/$�l�t�>PvD��<�-�i��!�^�`v:��K{*���_I�F2i���m�~��k�rj>�S��1N ���#+�CAۡ-z(X�� o)".���L���ۄ�����c]δ�P���;���-����  ���{���pPv����g�0"�\�?|�apV�qq�n�b�������XVb�ȇ��P.����+�)�Y�\"��y�R�U�+���A��Q*ev%|��p }᫭�����or��[֖j�rvHa�}7Z���=I�5�ǟ��I�q������Pƞ'����ձc^�����d�����mXo�ȫ�Zʮ�}��ʺ8��^�s-�S�*妔�ɺ6�ZB���5.ĥ��=mkkٰ
�ѸA��.]!T��z���F�]��)�0w FS�x1?'��zq#n(�2�:G����´/�}&D�o�[�1���,��^+g�}Ѡ/c�i������z�1�r$��4�k�޷�ǟ#F��$�sf �ˇb�8Ͼ�����g��%���MW��#���$H�}̖�j����k�Ʉ��޵&�TӬ��W�E �=�Vˌ�s�sEձ�w�15��c�wuܜ��BO�楍�1��Pq�<�tKs���G!�p���	�V�_f_ܮ1.�N�?��\8�5�+T�bZ����$mnF�s��0o�]6+�g�����Jw� K���?���N��&�d��4,q�瞜�y��Ay�˔�P�ϗ��vt�۹V�����Z���0EI3���Wr
:\<]>a�﷔/s[0��Z�
�|��ڡ���vWh ���w�׉��ۯ��ތ!�T/쵘�j%aD&�ifc�"�����v1
��tY��	 �JJ	�<D�jQ�͜q񙦐���-����p���Ju�K�#Nl� ɰ/n�h5v�"���B�L��&A�e�W�=?0r�x�@(z��5k��-�"�
k��ajHT�r�R� �C^�KS�{b�@�\�@�m����,�)M������BvK�K�����S��3mn��!&�����l�e0�|��89c���.K���e,����%��v��r�j�+_(�%?QK��]��)�I	�-��:�^\�J�7� ��JS��&���s+\��T��ʻS*�8Y��!���٘<���`�aVh��᫿b���A�x�ȳ�����)�ٺ?a�����cu�O�$��5�4�)2��$h~����x�V��������co��# ����Z�-0�6Y.���9]�h�{�g�m����Q���5�i
Du]���W�Y�ا�F���m�Cu�pT���ԁ�����is�x�e��N�8D��V��~t��I�	�r���S�Vף�;R���k<��>�w�(zh��+��9uM�Y���ShG����	� *.�@��&b�.���+i���8JЉ�ܮ%4��Vx�/������:��>�J�^���\G	#{�j���i�}��a��˚��a�½6G>��Xr� �+���xgX
>��w#�F���i��ӊ�?�΀9���G��{Y,�n�J�vv�3v*;~<�o�c�^��"̓rm��+��"c��R4%�����)[�(�F�=��B-��Ʀ�8�,Y�a�n��/��<�"i\�Ϲ�I�G|٥���C�Ċc޷�{��Ed(!�o�8|�}oNELy���4� ?�P�P]4���
lC�22�1ܤ������P�����si�����A���Ub�N��-{F�"&�ҐcIh��e�k�����L`:��TP�ފdk���2�/�Ի9��=ΐ�`$ky�_�j��iD��p�-)�d: �٢Y��\(�������{
��)�i	��p�5��l���.4*`��*�v:��fs���ι|VH�lT6�5'%B���j�]g6��%B2�3��h"��6�i���K[�ާ���W���2����L�&�JlM�e���Y�o�yC�M��ٱA*�}�r/昒��RV��u�f$;���������[�E��pz�#���!n&�����0ogCJ�I�0�X���J�B�sfu 
15�w_�y�@���\�8s���5KL�9��:
b�%Q)����!3��lW��P;��S��u͉�g�,,s�E2|�������c��ˣ>�ZWL�7�eLsF�.mo"�����C�m�/����X�a����@1c {_��{բŁf�L~*�E��nbv{v}<�Z���)f-�,ߛf9���lh���66С��5)u>M:�Lʣ�R	���>CWI���>߯�)c/��{�U����A�',�<��M�Z� B����l�M��B,�&�׌@}���Q��'퐰LrI���U�X��z���̴E�[S��?5���?b���B{!*Dhp��Od��!sU��旈� �8^��ph��7}��,;t[�>h������Ui8��&Re��Y���ܝ�����͎�v���߉L�î)9�8�;�M�I�(R�̟C�ԍŷ]�YkA�V��Iҹ@�g'����a��>(�H0P�(��ZM�zm�1�,=_��л�WY{d����_#�fJ���/��e�-T�F���i}�4a�4��`%;�L�ˬ��2U��@�k[1�V��^K�R,��6��!s�Wi��aۂ_oͲ�ᬚUr�7�; �i�.%���3���ɵ������1&���j�<�l|3��=G^�_�f0�*=���K����s��q6&{��G� �L���ơ)l�硑#F�g�������U��K�艖� ���>_��,C�\+2UQ����7]s�T/��	B���xttuB_aN�a{N6$Jꯪ�9p!������U�ԈA)���;�Cy��4w��<��gz�3�a`	��Ny�挡���vߡH��9�>���bVP`��|\���xzFJf�sV!QQ�ä���(E���S�F���E����H��/�}|:��Z��z.�Z�����夔��O
��"��)�����\,�e_��#�:�Ugh��ZI�e�/	�4�YM�2��%2.t���~�Y��J.�T�ƞ����'���$d:s%�����[���������m�W��8<��b�~&�T���"����*��c������/�C�i"����H��cC>����-x/�M���]�l�"���_����P��@k�!��)��^l�Q5aP�J)zd�����K�4Vh�?��!���Y���:^J.���;�@�_1|Y1�3�X���u>\Q�/;h 3#8I�Ӗ��:UJLEAý�����@�~���!����W<|%R����pSE��eHi�k�v:�e�.���`٢w�����.n*�Bw3;gve`Q�/��	ß�f�f�bt�����ڻ�Ȝ�쒒ӽ'�����·<�%�uBm`MZ\��BAy�3���*�Oз��]�{Y�i�7��+�N
�0��L]5�ר�ܘ���:PB�At�練�#�3���?		�|0s��Zpg&TғN�`C]#�[�G��iҥ���zqC�S�)Z��A�4@�d�$��nũ��l�f}RVd4e�Q�\
m����5�=誋T��e�vᨍ�K�0�ӷ7��o7��P|���yG��*��GsT�o�2o��А�V�ռ��.&�>g��_���bO-/$C)�3ߋ���D�Qfq�ހic�T�'{q���Z�Hy�o�ETƟ�8Q�:Ko�U���!�(v�"�C�nN]���p��uAy��>�#u��ek�aIt1p@����O|vf�μ)�~�a3����I����#qJ��]����5B���8�_9нcS�S�M0	��!?ԗp�D$��z��=+-P��n�T��2ٷ�m�Mݿa7
�t��!�9HQ4����=4��e��P�� ٠����Y��V����SӰ�!ga%;(1*U�;<���3��b�TY ��c]q��\��t\��f��m0d��T2�~2�i߻1ykIa�Xt
��!j��Kߏ�nY��~�'o^-.�������U��4��{�K�LD	��W�vV-�RĞ�c��pb1=����4���)�5l.�;��Hd�4O��r~�����>��`t��	Xy����Lك���7�~ѵ�� ժQj�/�-�<���Jo�������rx8��U@U����/gg��������v�_?�-F	:�}�k����	�a�wk3#{k�.pڅ͔�����kT@�H����w͑Եh߱�C!S����V��	��(_�{{����P�n��-���[�˙RK�'"?V�҅i֋�$6�>xɧ:-Z:�:a���_rs��iL����s��M��Q����{$����o4���1ke�7#c�����$bi-3����"Q1�4o�_��[�]K
Bug�*v��:K �pޔ��u6d�s�H�~з�| A\ݽu�;�\&�}�~y���SuT��k1�08��^K�WDK���>�̛d<�C��@��iƖn�&� �8�_����� >r�
��&�?�"$�;�(�gf��)�AN妽��|��c�BT1#|L�oI䒅D���e�,����F=ϲ�(��� _�����˖���L��.Mp@3���5î1��a#�g>�VC���	�f���g��Ӭ����t�o#�u.t��m3si(�1J�(���mS�,�)�ɳ� �Ws h�/a P�;⊳�&�J�_K��Zu��ٔ8��T��w��SRͬ+���͞�1�R4F䉫-`���>#�!�t��"5����_,���yP��P��շ�`�*,��25n�>�le4ǌ��)�ړ<�%��_E�N�.>���Hs?�r[; �E�O���r�E�����g'Ai1�����c���@χ�EXθ�jg��6'.��b0ݐ��nř3����e�>����#�*]��K����=���
��8�,	ܳE��&�T�X��6-�ǅS���TKz��؀1�3�z��m,�8���'&�ո�F�`�� 	��