XlxV64EB    88a9    1bf0q$�p\qZ�n�aM<�0Q��<z�l�W֫�?��F�
�x�t���,-k���-�%Sˁ�~ik������!�<�3�;��껇��橗����o��A�n���[��`��I2S�<�~H�g-���U���d���*�,��ӻ�O6�_�Å�)?�����DI����6�X��H�i�h4"��nI��y�I"c@^7v�=��;!8�K�P/�߃2������I��ј��+�5�6t����W��A�j��R$�eG�^�Y?�K~�+� ����Ш�X�P��{���r�S3�dxG)�����y�i0r~r,����_�AӘe��T�|�x�9=b?'��W��&N�w6����wN���aN�Wm�̸ʢw�[/���L��ND�ż�w���=1�%md�E`��H�CeC�k7K�#�
R�v`M�ʴ�xi|G������=�3l��p��1��V����z��q��Д��U��~�!�z�x����,���A��T�p�J�:h9�w-{��!������4X+Z`M�3_4��F�XsPdt J���ļ���4�)�+9���w�̢?�lC?��=���Y�m�K����8���{�+�g�p-@Yu�	q���0]�D�4��d�Թ��k��2�ܽk*y���`BZ��h3��P��%�UW���L)�/�/��&���tN������hcΜS���[�H��:�g�k�v�qӽd=P�����z����yab->�I^z�0P2�KN��G�5���9���^�,����*H��~Pb��v`AD��U�X!�`������Fm2�#?Ot����4	�l��*i���C:=Uu"+��IW�ޯF#v�������y*���i<@���ֱ�,���t��(����fU�s)�/X�(�O��?��@<�L���o*_�� \���(�-���q�ìi���5 �ڷ��1��wdURpVf.�OWB�)���g�z�6 k����$��H��m�4�"�Ac�=�u��[l�J=�
���q��W8��C��=×{;�C���"��Ũ�/y�����F���t�����&�N�9�2;���\|���v��'?
"��8[�9s���6�Ǿ��E����7��̖�H'�Ps}��
�4@+C�L�c��r���=P��jD+��$���FhK���P~c���[0�h�������*��� �E'�Ѻ>:ŀ�7e_T�	�r�Z���u8a?EȺ#l�Ԍz���{g�?;�F�QY��GqQ���Ȱ���!+��ϳn�Trø�������G�F����$��	��!���ȝ���,E<H+�0����AuЄMk�A�������e��;�3NP��V�1D-�OGQ�^6Ɉ���g�K�J��+��2���8a#�(�FMǵP�unBT獃1��l���e=���O�m���]YK��
����q4�.��={���H���Q�j`KV"9��o��iq���d!xT�DMK��㉾�e�����"B�+�˝��}�+�)y�9m�!�
滳���۷[�����c�K��0���L���$9�k�P�?�t���F;V>#sgC��B�V$�"����h���"km�s�g�e�u��e;-փU��9�p���o{�M5�<f���]1��Qf�SC77�-D����G]a7�@Ü�%\�6%��:av�kzn�����<=j<\I����,�I���n1i� ޅ�
��x�.�`�t�{�4s)Kp�ȥ��O�iQ�'l �;�
,�����Ep��g����"�����{�/(5&3oNy�;��	���J^�T�;4B���H��#9���ɫ�rN���\#�suF�í~��٬��R*�8#c��P���}zRG�@7�Ԇ������
܃3�x�fD�prG���:���9���S$���7_'7뺛"΃��9xgW��)O�/��ԭ�Z񓭌�O���6w�C2�2nb5w�p��_'�3Ũ�,w�3�������xπ�������ě����5@T�A���ێ�qx�{"u�ct�#�G(�R��g�/��Tcv�t>LUX)��.��kI�M6��wybp
�x!��"HG��BX��͵pI���T��.�P'[1�R��bp��W>`���(
gbe����ū�`��5x�.ۺ���T���V�nV �!"��Z�Z[4]n\����IN��"|%c��"&��R�0X�����ʏ���tr�� �� ޒV�d���7 �&��d5g�gBaOp�:/�o>�J���3:�E��P:N���%8�N��q�L���U�ӱvb�y���*�'u���$[��$s�q�*i�6�@S���/4$k\��'<.��eo�@U�Zq��o,�ɑ�0��OR��O��N��h��D��+g�k�y^Ȟ�a��Ygl?uN�p�ڣ���5( ��K̘�i��ͧ�{U�n��J��RX�S�{iR���9�l ��\��7�>��
�s�b��}0��i�"��#ԬI�5^z3� sr[����'Y��Ii6AR�Q�!�����T$W��'n9y�[e�]��"<�Va���Z/^?�����h6�l�O��(�_&%�{<<���I��T�qۥ�B��걦�h$��9�گ�g��b������1�M�	ط�з��&��7E|���@[��t|/	r���j��Ѱ99Lw�A�����QJz���P�sT��I�\�?�JMP�����K�ŕX}�:��
�>(�$�_����� �x��\k")�<i}���R�6�����U�?��m��H47c���R8qb_��\1��PS�X}һ�s����,y'�v�f.����������`��gB���r�Y��C�Э^T�ڝQ��pZc��F����cU
!MY�rY�R��C��>��a0 �~S�|ϴ��5&�k��1���{���<[���\�@����E��-����r'�5��i���Ol����<����H�Q�d�4f��>��</���E`2���/�w`�i/Z��is��h�*E%��EQ���m��Jg�3����?���o0���u=���uy�)$+dod�<�7���Zm@�[�~vQA�	�M��${)E��x�N����<�>���7L|��i~��|4�Zy�a���L��i��ց��9f4y��h_��Y<
~��nةu�˵��v.��B$>��̗�oZqh9\���
��C�[D�n����E���b�F�����ӳl�Z:Mn�V�"y�P� ��dV��g��vv�؜���uJ����ù8�w�]���t������ln�M�af��7����6@������+�C�����Qr�����ғ�d�(��S�h�:z�4LD��~N�z���s}�� �4�X ��szY�a�H����^r͂��:�*f�B)�W��4�iK�^�4b�/í��I��8���v�;����m�NQ��'=�*#g���8{J&���wB#��/A��9�������;���X|��ɨHnqό�[ ���>���v��ٶ�^̱�I�l�.y4�G6�c�?�n*������@Jx�� ��Q��-��lÇ�����<n���������Wc7�b����R-����k�ꣽ�תJ5sw'�����^�*3D	�XSB�?�"�E�"���<��xϓ5�
6�# �9�\�7|��l�E��f^ed��Q�����[ЩJ+kP�#K8�ٔ>�3�u�0w!�r�.,���R����H�*Vw7.D�������+�ω&}�m)M]a?�i0���z�Iv@;�v��=4�:�л&�A��ܷ�>����C�a�ygN �am}62W,�xh �c�T[N��`^�Ҳ��e�*E�C,������r��74�C.T��\e�Np���I��z�O]�L���3QHZU#��g��x^�N�)��/��~����]�����X1X^�7<Y�5�J��>X۩��QX�g��h���ῆ\�{���\̔�O�O�6ل�c��~�]��pb�06��Y`HiT���!���C�����^M�x��
B)���V`]��q����s�wDLsy���G��*ͽ�{hv���_�H��b��܌�!ɕv�%Tnh����6�
��f�ӶUlt�FR�`�����E��Yq�vV,��F@M����qa��Js��O�<翔('0��)�u�f�2�^��\�S��C�bN�o� ����<�Q�o[�>�2u5cSh�	 ���"��NYﱕK�;��D),r����z�H��7lir��C D__Ki@s�a�6�6��k�W>�M��q\���r�>^<��yɶ��&ZH�4N?��]}{��ߗ���tOX�=���+�����7���#�Ӛ�#�R:���p1:Or�T�-����D?��M6CO��a*v~T,�JU��o��+J���g2�:k�#�Q��}{�w�0�K8y/W���	ũ�LЄ3~��<��c?9��GC6����t�[�3��N��-�.qn,�TH��x�� �@��V�ִi(�({�~����A��ǜ�f8���3��[��U��5���&uY��Hx��a�1LQ��y���M�fPY���<;u?2h�bI","՚"�b����є���@�jR�Jn����[���������2��-�%�I�Ղp�)�f�Y��k{ŀ�ף�h(>�	,�]�ܕFV�q�"�m����d��~{b�ԃ�0.o)�%T���7y:�+*�D�\��M�}Ӿ��Ģ'�A��[��l�k���t����w�}g!�,�&�&i?�qn ]F�H�Oѹ��4��n_R�O�B��Dȇ0�����.����K��w1|�n�Pye��I5�ِ\�D�����<�!{4��y,�6�;���Z����\�j�5�.!w��z	A����wJ�X���"�4�./4tn�o�7=q�'�d�g�
F�)r�lL�:�2-G��@~�2Օ��ȉ�����R�$��.�'f;M��n=��ȁ�qn��Z!��c�K�܈����ö&���7��֝�D�+<��Uv�����P��qAJv�p,�V���,���L�z7��(�~n�*��HI�!|��[z�c�}�,��:;�p�,h_�>>���츭�u%��j���r[�S�	k:���w�ޖ�����.�b��3��\1P~�������qT@ҍ��q�W�Z��F���a{�n�Bt_]O)����:��9��R���r1�q�.+���s�D� �7*����&����5��gF���a����m-�D�{n�@��v�(��J1��0���2Cn�|����Uf��͡O w����67Q�٪�`�5�[R�WP�6k����n��>���Z'9f��3^���'�����u;�6?�OqGh����&�����;3�@�5i]Y:�^H�Ժ�7�!h��UF��3R�u����꾱1�'����D�O�&�_ۻ:�?ğ
�lU������Ȉ@6�DӍ�y6}�c���fx��b�!�_������&I��OJO�D?pI<�����,P_�-�3)���
�贱�9�«�CK�m7V�п��N�;')5�.8�)���?z�Bo�,Sk ,u�G��7���l���w߷ǒ��r�X����N�X�MV����p?5��5�	��"E���Aؿ?_0:��R$�����p���M����`����QT�#���Yd_\����=J7�z�� t�@���6����HU���<˯���a}���-W�
"]}&dr�C�&<,�d��FvΟ	�!n���pD�"�A}R�Z�;�o{��-xO��̘|n'���|��(��*�k�%���mİ#�R�\7@��t���w�I�YaGұ�:��=N�UW켥��a�G����u�J|��_�?�� �oas��&,����RP�Π�Y�����Y�Hc	F���\�a��}��a��Wͧ@����J:C�6b��Ɠ�QQ��'�C��nW�`��������G��Y�PV5�u{�������i�����3F�{��A{�z4��@X�W���􀜬�(-��,�ո�4�ј֖b��σ�.C+y�但��.�h�P譃�
�R��,v.�<��r�l��d�Ndoޙ�������Q�W+-ͺBdL󼧑�Y[�S��:u'+�]ǐ5� �����HG�ej�3�N���F^�)+�C�����`,�A�����Z���.ҿ~�'UH�T�r7�Ɖ#���\��v�3z�	���,�Q�z�]�hz$�柯��0 X�H���]�-�_����ye�@09i��~.L�e�+v��z��@ʅg�z��e�ax��ӧ��{�,�9��İä�b���͜��G(�)�h��]) ���F��o%1	h�E�Zb��ZDx�[y���9N3�s�T��`8��L"�a��&�rn9Z���R=�.�4mc.*��F��P&ؾ�)���=L�U*
4x"3����y�HN��dš��x���}O�e�j��1kV�/�K♕�����~N�������gy�G���p�U~~��xF"R��`�~�����_�HuJ��ė�!$�Y���Hc�_7�W�'vnI���஥�%��L��w?ZUs�~��7WFN8�+�7>��\
Ϛ*"7��.ɂ[����)��z���]��p7��? Η�����8�cN�P6��bK#��L�:ɫ�@���`��.����5u�I}?�g�O�">,���Mǔ^�D�!;E�����I��"��G|M�~Jǋ1{\�]�7:�aAp �&��<�@�`��.�وZ��UʽF��_+r�ͧ�(V�J� ���n}��l���ua%~~hh�x�N��q.8����߲��s��T��:�vT��2}2˟���h�ǆ-�b�4
c�I��ک:�~M=�W�(�D���٣�O���}d��Sr����uL�.!�]��-U�D�=��^�;�Qo� h�����bP