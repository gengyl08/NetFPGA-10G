XlxV64EB    163e     870�����:L���Ν�b�W�.DK~�\���T�Ѱ >��W�ӗ���a���w�po��z3.`�ڶ�E�'R2}�?�ꨏ'��L��a����Ҍw�{lk>�
y!�gk��3A)M��T]��wR�hx��_�uڹ��|4��=����I3��>ʾ\ܒ��Lh�r�����o��Q��'r�C/�s�n吱��0`z[���|���u]񃢔�.��v�d�r� ��^��E̢��~���ۣj�k�u_g�K�&�h�ny�v�E{ɉuyao�TGwB˪�Y(� ԃu�J�|���ʾ�=�Ǧ�ӹ�&�4�6���o䘕g1�d����R�K7������*��x|_���,���~�o�}��5�>㿟QO4ͥ��&�ѱj��5����R��grF�����~S�s
*z��lݖ��d�W�|!�w�R-�Q�!Cg��g��g�a@[��>�EV�ohڽ�{��G�шEJ����ꝟ�
 P����D4cxG���p��5���S[���=�'?�!�8�yʓޭpj�d>���MbY���Է7�_/[�YP���M�-�?}�53j8ƃ�6H K�)�V�i���m�7٫Ս�\�Qe[�2���0p��L˶�\M�+���Q�'K3ݐ:.��l�`=��ɻm��:{���bʼ2ՆkI�� �5�_�_9� ��(��L0�o��<��z��kk�΁u`�����߿_�^��M�@���;�`�{�����տ�Yw?�&�.�&�u���4�r�',&8]�Gs}�P�*U�I-�^��a�P���WuK!�
�����7�	��ή�g��c3���E��uM9��$m�r0C��5��'��:�!{%lDq��gaQL9M����	����͠�NG�h�;&�g�xWU��[:r.�)䒛B���K�\3p��e`0�N\�í�uyYۻ�/���q�H�Ky��Q�ɍ�a�ץE<t�� *��FO�)�#�&�es���.�̳���.���Tvٷe��i�����A���B``q��d@-�G3��%�l]j&p2em�����:$,�͆f��cz����`�4�%iT���(�x/�����-'��h�8��i|1�J�zC+�ռ���8=��������)>5�F�NEA���\M�5�K���G걻��{�b;�K~⛗>n$?mg�����md[��6���PX�Y��cBMg�<<ᙷ�(>0��X.}m��Ƨ����N�_���#����H���6P#�[�K�exǡ�M�<��>�T¦D�^�T`�"�aAv�J�����=~oY�5T�OO�zvϩ��h!b�{�)�E{L�ܰr)*]�Ȉ���>�eC0�i�A 6S,��r�K��^��ߔ�|W<'v2A �j^� ������P9ԒKT����&26 U3���ѭ�~���&]�sg��aFc	0���_�_<�0�|L��)�� uL\)O��p�l��9�U�*�R��/�ɂA�"���Z5T���}��jth�9���J}�G�n���Z���^�5.�܄�ݪ;����=@��h���f%*�&?�� ����;���\+��d}���7�$'��m��L\�����jB\�Zd���0�0�Z�.��D�k1A0�x��7N��:h��o޾HW���B.�L���gE��A�1��J��� ��������6�=�NߡtE��O�©�C��ݎƠA�M��(x����ML��Z�t^p��6"-ujrb��(¿����\��6!�O`�7��U㯥���wQ���T���<2�;��R�F�=>s�ts�i�X���Q��M?]�;ğ�rk�2r�W8F���\�#bM�"�5���PD��/��+�1�3����x���Q��H��}�3rιQ+��+�F�e�j�<��U��p��9��lQ���%�w�aO���w��4[���� z���8.���ցK��h�Q�������j�;��>�k]�oM�@Q_2f�O�uB�|�ë̡ꤺ��.����I/�h8�~u'�1_�و'_8�+Ow��H�=ⓙ��uvY�_�Ca�!��J��wN������B����-��6g���[�q9(��}����a�