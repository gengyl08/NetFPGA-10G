XlxV64EB    54b4     ff0�����h;��+t�a�q���R�f�m�a��z��E,�V�������QE+�c���&�
Z�ƁHPk�*�zs,?+��� [w}:0W��M�#���2xW�:�N��G3��Q��j�c�μ�㭘��D��'�P���z�k8*|U�z�����dws�hcvR[͠�4Kmٷ�`(GA@2���g�\��J~���hD����	���? ^��w�c�Y�q�>U�s�\ZVV��9���R7�V��Aj�F}D�q�* ?�\Kw��{��U<�]k���1!�j6�p�S>��Yo��)�w��%ab�`���jA�Y�(V��v�D���ٹ��65��B
�̕Be����#�����b]�XtE��1�uu�Pϴ���.Z��ֹ��Q1�\����T�<���Ʊp��-�yԫ<��N+X���	`ŋOc6!QH�� -R��OLWW�5u�M���-�*̇Zs{�D[��j���t��!ϟ����Y�
G�U*�ǇѨ䢇:��֢���e֦����[�x.������ѯ�n�	�p�ן�`�z��/�@��Y"l�r[�M;RQ����ge�i�$�p����q=B�����+�a�k��G5�*����S�ڳ�-���z�/eY�YY�ҢSôUIH����l n�C�Dk�}!��=�m���k�.��?fd	��q1o7�U�@��\(�������g$=����r��K���@�u�UЃ��k��*���BO,�@��'��Jڑ���<5����n��U�6j�RЭ�	K���u�TeC�Ww��ԧ�HI\��K��MΤ}c��� �-l��ۅIwz��-$���|T��=�L/n�e���^
>�o����&/� u��n�s��6g�1�^��+q����;D>hB�bYZ�Z�h#a����*w���ҵ ���oi.��ɥ�8�@�Y��JU-WeBlؼ�Dv��e�v���fNF��/�ku��2�J>'"�+B��]�U,�5�7=��L,'0���S�%�ug��Nx@�a��U��Wux:0��ϲa�,~�Ռ�rS=��J���E������'���q>b�:گ�FD�]F"�`�^�2=39�E<����b!A���}�=�!�\
�-�L\�E�<�����Gю\�y��bƗU&�1�A�-`l��0����б�5�;?^��]̏��M7v�D	#VX�EK��4.����A7�+���C�`���։9���e��Qݷ�ۓ�\ӝS|�,�z�%������S��T�eP�y�S�&H�`Q(�R4'�{�Z$��?�r+yy� �Nӻ��j@������]Iy��7���`��?>������=3=�|(�;hb���_�����a�_��P�Ď���zy�.�mi)�)~7,+S]��U(b!5b��Q�*���˱)}erdp�_��1��<$R�l�j���T������P�J����m��ʄ���dL}ȱ�ue ;�8�Dr44ԵH� C�,�_�9ǽ��Pnj"��K'Mb�l��@�����\����DZ�r���v��E��Hb&��D��jҩb}�8���-�If�˹ȼ�d�˾>7��7�pp�8�-=��|I��.P5i�L��y��-��\�f���'''-�~Mp�쾘t@�q���N�"��\�ѸJ	���_�[�py����+�:���kb�rX�$y��O���M<C�h����M��a�����J.#��ՠ�xc%�M�4�\C�9����ЇۉK-�^,�G� d��X�n�� É3h���f���$3,�����o�8��b��,����c�.Yײ%[�;����L��x,�Ȥ���vk�Ż\��0B=!Q��$m)��3zba����6iR�qpRأ��P����6e�X����ު=? ;ݕtF_��d�8�Ի-H�c�(��j^�Y�`�����o�ex?%�?>����L��n�/�L�K�nʭ��3�![f�Tר"P�q��T/�/��%`�jm AڲEk�ҁ���>h��� x���e}۳L��Ԁ��Lp��M�Com�7|�� Ǯ��9�0	����"�B\&�a�__c_�������5]���7H��V�w��D~|�r�\H�-����gmpb�9�kh��U��$������.X�A�Q�;rv��t�as�;�UT4D�{�����IW�g��v�<��WXOu7g{��0!
o��$@�4���Dk��{_�d��_�_�/S�d�:iZ	�c�9��%^�_�ۦ�Tagwh��_1w��J����f�4�0c��h��ٰ˵E>/M��2}�Wk'��s���rM�&�g�g%8�O�sw�b^ث�X`n3Px=O8�Ĺ �k��$�^�d�mi<���ͤ\�ئ�ξ�Q<
ߢ�!u�� k��x|R
�*40����Q��T4E�H��ݬq�nx�7:%ּ��,�T���2Y5�AC@��0����aF�qF�pz�U��7��L��ݗ����9����d�DџL��y�B�D
Y�?�C���_!�Rj�ߒG��n�xX놪v�*���ڜ6�Q*(�1`�٤8A��)ߧt�Y���?N�f�ʲ`�'4X��}(%��U�IWl��(su�x'+�CQ�Tk�=dV���mF�Ag���	FY�}D�k�8'Ӄ��JPwf�<r�_�e ��8bw�{JK�҂���si�U���%AV����EsF�rCj�Cb����tt0�̝�-��	SA�+�nß���f�N#uv����4���X����Ɉ��/�Mp�f�ou�U�'�ڂ@Kb�&�4]������u"s�ً�/�+V0!�4�/p��&	����r��A�V�͚@��v�܋�j��t%b2�mI57����a��ÝNo�5H�uԡ�=e.�c��p-Eu0��Cw�\aG+�߰W�	v���	-Ѕ��0ʱVkT�y���zh�3���6;��c�M�t���c:�K2�6DAж����o��d�E��Y1��L��u�z3��Y.a�r���Li�,2Z�~���C��"��S
q2F7��)�%-�+Kg*� Z%V�:9�%�B�T[&��*=6��?� #��m����2�8������J-��j�:����6���p9���`w!�x' tYv~��%�P?LI|�j:��j�u��6��C����e��)��� ?�NNsxI��P���+1H?�9�yY"s(�g�Z�.-h�r�j__E�J�N��|Qńd6�j�2���Diqav�a�4��]���}�F���ր6c׫�I��|�G�+.��JI�&�KW�=��P�T����b���
�j�8v>����T�4/p���@M:�.���ÚrXN'E1o�Ve�Z��y��1�X2��E��Ec`t6��i�ѝԷ�{�&�͂BQA$	��n��1�c�oN����˴��ݰD��4�,'�����N�q��t�0�֖�Ԭ��:��.b����0��	�� ��tz�tx�>]'h�r<�F�X��}�.�7�H.M݆�6>����P+t!�����Rw��%����o4I�BKa.w�A������
�Qa���v ��%��z�3B\�	}&I��x���8aDG��~�וE)�5�}��A�r��\mѰ @�����yS>�����a���~���A�BK�S�E�!� ͭ���nx]ܞ{H����4�X�H���s�|E��cCx����ǅ뮐���:`jX	5��o_�������$Bx��5���d=v�+)�D����AҘ����
�g�=��>�5�-���G���(�+�&����߆ޝ�;��k7���9�J�0�h���6
�=�	c�6��NY���c��Lf,��w�E�_��a�-Y�3�ט��ڷ�Wc���=�DL�HεZ��qdC��d."���xϸU��br�Ld��K&�|Dɗ$:6�w"+�0V���h ;��󍇈��u�&$<�J��A /�^�
�ۼ����j�]ڗ���I&���=��������1�Sߛ