XlxV64EB    1dfe     9f0������*dxu#¥�x?�%��V	�&��;:�	�b�q+c�h�xr�����6�(�u��r5�E{-_��nW<�׽�+Ǳ�)�����6B�����t�b�[�V���R���4)|�K��$�d��I��K3��wAH��+��q�:�e=�i�s���?�,�泏)=�sn	���8}JȂQ��nXj/����~*<gP�]�b���K0���\��+$-��,��׮o�PFyȩ�qr��b�A.���d2Q��[`�=��,�Y�������e�J��s���f�9��w�GCc�CZ%��H�d-���gO���[}��Q��������B1򼙃��	�	����������U�v�"� ��g5&��֣
�EnZ�m�W3�g��מ�,�m���t]��9�olN�@İDhVg_i�`��l�
f`�������g\�֒��<�EŽ��U3P���i�Ĕ@Cm�U6�cS�#u��3��J�"����|�?ah{��ֺ�'�ݞ�`0��_��̝�]�����R@w�i�� ƺ8?���^Y����u]~f�I8����U�]I ql�9~qNb �s�)is�ZᔌM_v�������d��%�㋎eG�N�b��Q��$�9-���?���F���K#YR��L�8�_��|�}�؇(.t�1MX�c�֨�n�R���u5��pVƹ�F0r.�,��L@�mxʧ� �y��G(Y!e��ΌGn~�V�� �(����|�ϕ����D�<;�F�|L���ལ3)?�4gS]ѷ�J��k������0�,2!���{*Y��h}�׫GI���v�Z�Al������~S�3bU���c�WL��H�϶"��W=� d�ʹ��ɫ,�B*�K��8<P�Q���y��v5I�eğ6���x�_5a�.�M/�:����2c��V4As��R��������h�dt�w-MƯ��ʲط��8c>L��@�".�L%��A2T�3�c]" �ϳ#9�~�R�z�p+��7��w.�U]^c��
��0����ڥU�X�H'~ZHj�tUЎy�B�#���-��lΉ�A�Q���'ۧ�́�	p�X�Zt�Bqx�G�:��qn��z�@�8��9��YՉߞ��ܾ:v11q:ğz��P��VG�_����㩳]/q�!r��c~򘽙�7����YעE-\Zm�k�U��6���m�������C�2Zݦ�A����DZuX�
w;�:��=߅��;@8R9A|p��i��i��v{�s�9���QR�.X�;�D�S���������o1g��Zv�;PX��1ܛ�dg�"~oD�w������M��H�f�*Y��	�ȟf�D�R�YIHd�k$�&�6�A�0&��+���<�l������v�p���prﮞ����T}����(���
U'j���T]��*�lV�00�Cc�5��^�����M~.��w��QM�.�mB�E��$��� 
�?�0�qI����d����h���qV�YO
r��^��xEo�+��8�������YrƈS�x����Abtj�@eNc�ĝA��>|P)��>tj��m��d�\@]8���qp�`)�9N�Eq9aИH5�A�S&�7��ʾ#/B7y<t!�L}? |xGbn�I%��Q�[���;Χ8��_D�Oh$��OTs�ט��iԛ#�2��$�7�|1@o	��	�-9�C��W��K�p.���!���w�/Jz4%���dʢѡO�]��>������_�����SCFoG�x�[^M�M�ة���w?�n�1��]��O����ZCC����Dk�t$�o��V������Q����
|.��*�H��1d3�z�R �)����n�] ~a%g,2��sf���8Y�t!+�	_m�
s���ˋ�|߅"��!�;)����xS��p����4�z���7%S�"Zo����9���yN�bGj��m�9e�E��sm^K�y�+[�Il�CŔ���ˊz�N�6�ۛo�������L��ߔ��=�U���2U`�3�(�M��Q#6�I�	���,�W�Jx_k�9�ߙ+�Ug�"�4�Hn6�B̰��j+`ęWz�C�7�8](쉺���9���)��;i��7�e0_n[�D��>ӆ�1$����:}�'��m��AU���y��\����� ��GF�Fkn��?��8���@��Q���չo}"`ž��Q��3�?Pf�z���f����m��Ք*Ɏ��53������eO�`�@�[�._:�2��R8n����-��&Ix�£ݥJ3.��1���>�#It�oA�4���1��%Uj��~>�9U\>-0�!��/��K$>"h����Bep�N�q_i�6��* �.YlA=��}D����ma%�'�1�|}"��T�k�NLG����^��|U~�۝b�7$~�>�%9[ih�/�4�0��AFPq�fx��p
j����2"$h_�����JW�����