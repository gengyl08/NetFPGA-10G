XlxV64EB    23e1     b50�"Tz�*x�f�ͨ�h�w+$Lw#���?��y��[R(]��|�c`�1��Wt�
�x;rǌ��Qe^|���^x�u�N�E�����<s���y������׳���5�g�Ψ�u�rU�PXM��.�K���l���(������F"�"}h[���(�wk�q�4�𱗆n_�.cJ$��6B���	:f�G�R�?�����!�4����i�ӜE��H�2�(��Rm08�Rj����CHd�J7@<c��#?�2a��=�J/i�W䞳ǝ��z�a���1c��Y�)[���0*C\-ɋ�߾Aq�}�OI3~�v9��[ʽ.��/���
ݬ��N���G���%���v	��M5���X/I�P�[� k���������T&a�^/[h���1n��C��i������n�~����8��y�cIxȞ�v�ν,�u{kU8t�/�&�P�{KyX˃��)=7i��H�^�q��2Dp�I���bt9���dr�	�#�N�����0 �BZ�q���^���M��"V���}a}%;#I�ʝ�Ԁɡ�ӹ��`(�U�P�rzW�P��g����ӻ��U��JU ��=��ntF���RB"��i�<j������7���s�/�o���4!n���F������޴�v*#�M%�� ���vF���l�qAWV���h`��u�T��[;� E��<M��e��.�8������m����,3����uL]E6��v�W<2��S�27M s��t����%VC��2�����!C����H�؆<�V,�|M��k�z#&�zD�q�/V��</<�i%J��-�r� ��0�xf��b��E�SU�}>h���H�D�O{��gñ^�L��I�r�k;{�M��1T0�d�
���=��DL!�(.؎�s��*p��LB���Ց-�ynh����%'���Ol�LW�f��Sj��/&*�M� ;F�V���y���zei��!�C�<'�9'�Y4x��w��X&V
7����7P�+,!���u�y�]��૕��ŕH"ƹ����(n��[s���� JgB�`��lŦ�V�x���-�2�k�<bu�D��T�T��H�L�9���2�2�no��B�P�M�ċ�S����\�s���2#r�����5����m{
�L�r�i��y�ΊL�\��������Ξ�j(�[~̱�ԓ���*����k�{S�e[�hU�ZA$�"��Ԏ�wx�`q�1�3:�I�Ӽ»�y��fUE���?���WA�&�ƨ<�pW���tN������8�p�C���㜨��{�j'�-_#���P�"��o̓�.Nr	=�`��n&q��y�DU^���G�麘�2S�'���nv��%t"lz�����`����c*MX�z1��%�<w�l�����Îq򥡫�0V�rw���PHauW.,q�!�Q�T�M)�"z/�ɭ��rW�1�nR��&?҅��ȿ��;O����U
7S\��FsL��,��)�ab@���q�U��2vI���.�������L�M��8s9����c����g� jؑ�Y��Y�I@ET7���{'3�{mI�'� &kR��s�v��������
��L�	�Q+r�p��"���מ]jsP)ߎ�%���Wx�6�J�1X�j�2�h΄�
���JH�g��	�~�����)1#���4Њ3�Z?�K����sGx5�y�����-N���Q�C,E�f��v0@V�*��g�5����<+cEh�mXް�����h
����"��~���w�z6��;��˸n���R
<.�\�����U���A�jQ� ��C!���YO��� <21��"����P�b����{DUy:Vn�d��rPz8'ȥ��g�+��u��y��O`-�n��`�	D�����~�5�"�F� �C="�nA����8���ې��f��P��#��6�?� p�4�$��_)�j�ߴ�E2�AjZ�r������~k��dn$p�_)�}z��2�g�d����cʫ1�M=�@������LF��W��3~fj �����[�m��MCJ�[7p�	�G��2%�p���:�T�)�
��څ��[����:���pR)�a,�Q-�q)i���V�S�3^*��8H�`�;�/%����C��ԗ�"\�7FX�5!~2���@ t%��㗍?Km]&��~7�67�B���<Ƨ�H��G�Cw~�{q^*q�Ogf� ��G��;Xy����W�ђNG#L�N}[��G&.��5(�1�L`6���hM�;�ryDܛ08M��K9�y�{�L��k�/))�+ ���'5�@��v���T'評<�R�m|ݐ�#�#,����&;FP,ʒ��/�([;�@��6Q��fRaG}�!�w4=}J� ǃ7*ӗRK�R�!֑� �� A�;���vEPU���JP/�����w?^�F�4�Y�,T��T���u�=`�T8HYo�&Z�Y��(2�eT̼����_Ӌ�_��g�"��Moq��2����$�����ĘJ> 
U�pyQ�&-�H�ȨNJC�wv�y��c8�t��bF�_V>�d��m^}��ti��ߡ�Ztߗ-5	�U�	&8���հ~����~�^B�)��I�i���n+a�U�SY5fv��AԸ�D��'�'[� 0��[����.f�n(��=֒�o����p����� ��������[��gLo.�6��C
y�;�k��av���|iM�QХ�c�}4i.�Q���]tqF�n�燥�]�x i'r�h��ݡI��s�]C[�b^�-D�^&>���g���?3