XlxV64EB    56b5    14a09B�%�=z@�<o�~�\5����k��V�S�q��[� x���caɁ�|�i%�VVx|�����W��_?U��Mkv�t�����Q�6��vF��2C�-_��t�%��'t9�vI(*iW�S�T%��h�n���5yӮ�\����m��;����"ZU��[���[�z��'d�r�wu�x}��[o�c�����h�o	�)g/0�����B�΂N��V�\!��<�Hʧ�hVN>�?J	E�1׶"	��R�����gn�4��D#�A2�c�H��&׻���h���D��#v2�!,���`�ۋ49Ю��۫���e�n�ߔ	�f�(��Ɋ�7�m�"��*���������hϵ�nx�,�������ty}%|d���t��g������v�x�7�/e[��⊣�_j��֤\BLk^u?��}!�s�!�[�V����&�X��a;͡CA����.<��p1eW���0M0�7�hk;>x�������w��G��۲��sU�R�Y�a>F�jG �Ll��1�>#wh=�&ǼE�R�B;$�IJ�v���{�N0-	8� �0�x�/�u�k\㐼-J�
��`j5��.j�"��|΀��x�Hp�q�]����R&]�v�tδ[1*��m@��>2	�%�Uǻ�VV�'�BaUO�Hj���z�]-���m Q�$�>q)��礂��T"u�G���%�a�]B�<��=�S�e�
�6�7��,�*sn�\1��	��-e����`���x�BB��)��|;�[����m�E���=�56Q5�`D:��)��J��n�J�b��'K7H��R����yq�"p��:�9�H���B^�s��C�M�㭩B*��X$�K~J�'t)ٔo���/���P��N�udP
VT�B��U��pk���~ض��ƛ�o]�m���/�WfӞ��w�5��lt�lW�b�����|��tsZ�X���z^N�w��̶d
����\א�A�U����(�D�R[ ����ZwA��hF��h��{����������O��m s������;�mA��֡�Y��+v�ip�"4N_��4|@.:j#;ϩx��gU��L����Ee���Bĸ�\=�+��������ׄ�^�?��q�^|�a����V��D��Z0}�~��^;5�x�0l �ɟ�֯�Μ@�5މt�i��כ�Aߛ��gga|�jS��N�i+6�o~
O�S�l��5"��S�1泮�5{���҉(�D��V�p6�-� �d�@ܩ�o�W�G�.?���- ��=Ѡ)f�I�(��qcu�=M����RT^�oSΩ}��z.�`$�0�c�R><��9�ݐ! % ��׵D, ���L����Е��y��*j��V?�qfCK?�-N4b���5rx�^�J��c}jS+� �~�w�B��p�U������ #��:����&��8�}�^��F�(��O0I!���b~�י���� ���8������%��� ���LC"c/U��^��3md(�;Xj�}�i���ڹҬWA*�[4w9N���s�Ls�߷g< ����l���b����ט�,�y�u�S�����A��^�|u*��Ov�4�+@ì�;��4��g�#��=�aie)I�E���A���]q�<�[�*n^e�%!+%&�ǭ����-�8��	s�����z��HsE�� b���$z���3�e��ƻa'b������Ф� �����[QL#�/��?~��ٗ�(M)��B�d�� 9�R���JJdU�����gz��p8xC��#]w��tމ�g��#r�7���r� ����f2��%���I9Q>Wc�?���}��\~&���J�!&��c~�Z�X��n�{Yv�G!��=�_j+e��Ƽ�����qC@U�F��da� ���e�	*�Q�V$��B�6�q�Yd,N�e�'�_�娔��o�������t+¨~�t0�E�yʵ���:���HX�P���3n�]#�W6f2�JeC"�ã����7��n)|Np-
 B�r>GP��/@kt���C�c
S �=�����v���|Tۃ>؄�^�
���YR�莖:{yh �0S֬2���x���f|+����	CS.Gp�����k�6�N�$��Tk(Vu[�_"W�p�ȟF�/Kh@�V��A�G2fŸ|�21V�qh����i3<>'7�m�/ђ���bN��R-�����7��6M0`����K�S2T��_�F�"����p�3�mS�G���^m��I���Hqt/Z�	�U��c��,�Εq���s}lQ��+s(X^�L����<Z��+T�ښ3�4B�:����;���©��͟|�Px[Y_ыH�rwr�'D����j3O��(�9㉲������a����ž��|]v)�ŖB�����Q������\�K�T��<�сb�'X\�����d�eN�wE��/2��.��&3��b��48���[ ��_�t�s�p�_�H���p�z�<k���%�70� ��D/^�������v_�����Y�}�C7[g��ʐ���/�UF"#�ϛ5B�p�M�G a����Ϝ�ݴ���I��1lU�˂�p�rx��~dL��4�N۸���*�f:p�K�!BH�oE�m�U@ �H�60�,�,L�K�܈Df�e�>F=ZS�C��$ŏ�P�
3��P���~�*7�7������i;dd���4��p�%�� ]�}��j�θs�:�ZG{`Ιy�G�������]A���ʷE�_/?&��f��>��Y�������2�n(i���S��;�n����%
(�Ֆ�0���h�R����O�Hp+(�1�\7��( WK$5�:~�7� �WU�q3��z��`��s@�?����G�ʿ"Y�jz��?+�J�!6��I-����%�����eMH���h��{{��#z��fC:�z�	�������ʛ3�e6�$rgUzI�/?a�Uv;��P?� �'_��Y�XJ��m�d�S��	{|=���-�|:CE�fL�*_F���}�����_}M2�u���$��f�w���.Y�cY�M����ڱX�ɽ���Vy���Q���� ۛ�4�i��V/��y�҅�����p�t,�����")�GS�U�%w�`�mU��꼮N��8�1��)g��'e����C�2p���lg�&�ZjOy��Z�;H�M��Y���Η`�C1o@�������Ea5ƳW^�q8�'K�?~�`�N�����-e@�~��诣`�t�p���-�p4�M��c���ǉk���}߶q�n!E-�6�.S�?�_���gX$��L{2�\�O�wO%���.�w��F+ cro�mm��M�:��N���_\����/(HM�b��"K/����mJ�.-A��H�.���NplD��Ҏ��:|	Xt�ui��7|�(�]��U���p��������߬~?���?�l�@���H� k|�\e0F���j�r��8`@�۠�]jA��7��h����HO�qif=����X�@�!����4腌*����p��Ʋ(ys2��o������)�g�}��V�؛�^m�zKZ���I�k�tW�#��D!� ��|���T��glg!0^){�n��:�b �d�rdQ|���sz>������6�e:��k~��.�e�/�\=�UBo�����W���1�3�~�AO�`���H|\X���c/�U��R���P����d*��6O���کjZ�����C�e��&�S�F�!�LYxI2A���f��p�>=��m�i�a��W+��BN:b�9"7o��ʪ� l�N�g�Y�P�����)9�Ʉ"|f2�s��]U�X��w�� ��Ц��n�XBQWCH�ގPIV��"���#���S����?�|&�1�3�G��zJPa>�����k$�uw[�9)���ԁ�^ݮƿ	�4�؋׃NqC����KҨ�̘�%]	w[�J�UӾ-GA2�>L	�?+��d$��ߝ�~䈮RN�9�;�x�p�2l^TbKwz\mC�ڍwOaR����Wқ�9(�ڳ��Yj��枆U���]W�������S���\܃(�z��*U�Gﬖ`o�$����'b��'��wX�Jߙ"���	�-��� \�TsK�$��B�����߆�1`h��ͽ�;´�0[eN~6v4�X]�\����+�b2��>��8x�7�½�BM>ݲ�D�T�yk>���lP��Xc\�C/��A�}ހt�Q$g�+MDj��Pa$�{~��A�?e�7C��V�).�a=�.wޫ>@�=�|�q6��	��o�l��1K�����͝HDI�xTe��^��[3��$q�o��v�����Wg�~ѷ��e�Io�^fw�w�֪�r���`��I?��b�m%�(�m�u�o��(��=Inw�z1�!�$�'�־�K�D�!��;9���!P�BI�-Id�+������N�.
)�}<�8���Jw2����,=$C���[3�3A{�����D��\40.Z.�@�Q����ćV	�1cR$�׉�*�.�J�[�.�vƯܦ��~YҮgu�4�W�Y��5�86��I:/S�b&1�3m��^��$2�Yd��i�ݸü7!�E�$��Xt��:j}~�?��Ҽe8���;�nǃv��r��󳻷�?��B�ࣺF=P'q�[T}�t_žk�,Km���|�P����@��_H����IY�r��9Ƈ�b�J���6��;��0WPI����
q2�����L�'B�)�A7D3}H_R�[C�tjg,zX��/��1p���u��9vRZ��¯r5�%��qr��n^Պ	cW�C	�r��Bԋ��[����IQ|\=kl�l��`��'��M�|j�dׯ�Z�9�r�"�(ع�&��:�K�l�v�Ӑ�pв����<�Q�ܮP^~��;��=�����*/ ��_G����O	
� �D�]eTՄ�b�j�S��(�_��B����#�ò�������A��{��(��ME�IW&L~�FY��ވ�76��=�{���_��M�- �sŹq���Of�p�`�@�B�)T��\�r���HS-�$��o��؉;	��>��J�K����JX���J=��O�W�:9�H�Q�c�.t�T��{<bԝ��-�C��͞��K�N