XlxV64EB    25d9     aa0QEY��rڍ�����lf&���c\�W����t\�ʪC�n�ƈi�xԮ�H7_t6윣+�����@��~O�L�Tc�j�j&L[���!J�EmⲂa�b��g��gJ��af��[�����Y)8��1�ҨK�wcw63�G�V�fP|:�&Pp�yPJ�PFVK���񮭌�}_��'�)����� �o�Z���ِefv���X6�yc�J5n��2~	��-D�8_*������vH\�J��댵�����ͬ�"GO�sr_�@�,�}�ck����+���(�M��D�v��6 �������h�ԙ��m���ZLя�g���*^�Dǅ��3�v�%����2�+Ƥa������UK}?�Hq��� �Q<|�?���?�bT����T��GIVf~�l�i�;RM#��� �|5��
�?��υ�g��q:�-֘�}D�?<�i�D��?1���d��#Ű��mhb1���m Z`��_yV���5ڢGG��f����PY��:��@�K[��sA�3:ƕ�Z�p��a�C� �f$���Bht�P(ܗ�F���p��^F����uR�w�y���m�����ᓂ�%���0x��T��-ܮ|&ϼ��<�;�"CE"4��dQ��e�C?�N��M���tA�{�^#M�t�nY��ۿ�aj'e���9c#�^u���bɇ�|(/.:v�W�I��|
ﶅ4�Mc�b�!���xT� ֦�Rx��wN�a�.�u�q�R���AUE��C�'��.��8.?��B63ʦ^�-��[����E\���&��D��C�H�~�8``���1����f���o�~�.yn������В{�����0H�sn����V1v�0(j�G[��F`��d2`�����-,D�'4�� ��}k���QQ��Ś+	���+��� ���N]�Me���H��:e�éNa���s*�i[7cӐQxG\�y��-�I_�W|l�m�@�*����`}��L��QZ*
�;��t��"گ�f���g��`�����T��U˱W4�����U%
�<k�>�`�4�4�I�����<�^�#��P�
.��D@�|K�a��2�:෋�og5�:=��Ό��"����_7f����ot�Xԗge�-�Ez��~��D�p�+0F����a�E�#�PcuG��v*�sadXXr�41�'c���7}�l`х��0g�)�ѝ
5�3$���&E���¼wL�[�G�N�w��v��h��e�r���Q��]鏫�32/�9���.H��Y���̾��Ю���U ���O����S���U�ܻdX�7�m�;�2'yc���J��//aJ�Ym@��Ὁq�!��dz����C�vws�2><ܡp�%���9��W�	9��R���i���F��$z[\S+Pz$B/�p���H�V�-n���n�PӌL1CF��B�����[;f<��^&��|m0I��􅶗��W�w���PgW��C�k_��c��HSԂDAM�Z�˭$���&ӡl,и���e%w"�)I	1�5,��˓��:)X����.�[����i�ij�7�3T�4�!9� 	'H���n���Y�׉g�>��Bx�=T�]��Q�&g�R)w>A%��ѱ�mr�WӒ����z�W٧w�V�=�]�y�
�N_i�9�_�^�q�P�9\���k#�I�L��3GG����B2�e�BR��a��]=Ջ�"J�_*~���#9�K�k��+f���D�i�$d4��p��40��Z���:1��@œ�*ôh�����s�K����	�
Ŭ#��k���Zs(�����=����2R��7q�lGvr#�9��� ������#���|P@�5`#���ͯ*��0Q��̭X��ۓ��x���M�QM�"��I�q���|.������},
������If��u����UNz���p�
�u�B��|V�f\���1Wa.�ƀ�}*vl�s<b��Z#��:�����k$��������G�*��&|H1���|Lw���U'S��.�dc8A�>3I	}�b�;!�}�N�]`4:�п�.}�e͂(fK�x8M������|��|T��I@�E��b�V����e����$��:���'�%�m��ը�n N�ǌ�4o����7�T�Ɠ:�R��=�8�x&�Mw����t�)���z6�:ڤ��	�M6-i�I�Ng��*�NIPr�̳1!�$M�Q�}T�PF���T��d�	n�^Rt�!�A�[CO�*����W���Cj����C�e4�c���{2�q��}�8�/ʙ�E����)d<�e�O���-�D��V�Y4��H�1�	:���n]Y\l�fڌ���˱�R������y����ٽ�mA����D��i˼��x���υ�Zot�#��`�|^;ܺ�ם���B�,�e����d �~R�=�	b�ņ|��0%	Q�I6���q�����;���ef�3�?PUl�� 5#m��5���I�@�|��C`k��q�E��5MI��h��G4S�����d�3ws*�����I/x$ [�,��>o\΂Lq�����OS��
D�PEڦN2�_�	lv�,3�\8@YjZ-�o�NfG�Y:��t�w�re�H�H�#nQ2a�1��E.OG{� �Lwݞ-��"pM5��FВxx���Qp�0�