XlxV64EB    4c5a    1470�)����`*�
�g.ݜXuV~S?[��ڽ�6�f�mF����<��A�'B�$Z��R��#��O�`Z^v /�8Qjh��[�����I������/kE��7��'4E��2�Ӊ�挫�Ә���o�:g�����7��H�;o�֫�z ����W���R���������VJ'4��Ԅ9�Ut���ͷ�0��d�����j� ���d�=	@Y�b�%��	4�d��GR�5=��B�<� ��&������uS�u�²Uϵ�ތd��N~�"����V����&hF'����)@@�l8�s�i��\ݴ��x �������]f<Z�3�e	� '4=�6���Tcr����Ƚ�ZB�ըd��GyƵ���	����[6Q\~����ߌ{�V��j�q��H荷�����oR�4�Ǥ��~���j���Og7�zT�-�`��2*�Pk��'����5a�}�)�G�b��IUGdm��v��y;pǹ���E-�W���I^\e��6�N��
4�y.m�8��2e��5�/����U)D���<,�E9�X�D�"�f������u#���u޶�q̜�s�<���1�?uw\�_=�}eW'�-�s�����1�ǌ�	�
�;!m�D�T}����p	�ܸ����0�Md:���B���@2�q�eĽ�S�x&v������}��"�aFh����F����G]+;(�����9[�nѿ��,{3�m�fS׈]��f��Gk2�������'�"��^��|in��M��	�I$�C��ǁ鵌_(n6�A ��K3[��ΰ*�h)_��w�H�,��Mx,��z�w�9��6�G�V3N�U� C�Ѳv��[�U����t�3��--[cF����l��WF��>y�sh�a�囚=��N(!{O]_�KN!Ra^2���{n�eP�6(�͐K�f����/G�٦_�W��$b�[��魤N�7���n8S?[n�/��EP�VB�G^�W��
���g$r{,�A������
׭D�����y�v)�b���ւC��8-x�/��W���x�h��12S��i�)�(nV#�*�ܱ��|F@JO��K�ڀ���T��=���l��M�U֜�h�c��_���HW�����\9r��5��Qt��[�
۴�7�h�I)e��"p����oBi��j���%�@�}ܩ o̿p���/*C��9?�i���xG$L�%F+��~�x�UҼf���רa���oA1�.�~���]SFF�EH�(@����@	d��P
	�S��ڶ��qREce�	����-��V��uQ�G�k��pu�þ}�8|%���WY�66o�AO*:|IN�1�v����pVC�M׈ah�%rcUa�9��H���h�E���r�X�xt�  F�C�? K�owo	Ό����	�/�GA��-�Y-.b��tK[e�&�K��}�+���.������K��-��P=�0��h��!��}���-Ec���K}1���n���!n\۫���^��\�Xw�2
E�*C��"���ίjZE#4|0�H�0%�0�#،)>��I(�ݨ/�[]�ڟMh��hI�P�qn�^Z��ax��6���^��Ǧ��5.���e��\"���Վ�'���	�p��v��lQ�O Kr�A$X�Nt<��Mю����iuQ`�����u2�]X"������u��Tn�যi��8��~Q/7��yqAIO�n��\#�q�+��q�pմW�Kz�`��X7(V*:�r����W�D��Y:B� ���?��b |�
[�"_� �_�p�[FS�;fwd��:#l��=�bB������nLӕЏV��iɞ,���Ur����!�:�W�c9ܹ/j]l_��GLM�ZW�p:_h�R�0;�	J�M>����7�8��l��� ��Nw���w_Hʱ������Ѽ=�Lu�wTqܸy���`>��p�ѮO͘�?��rsa4���\�d�u :#�5��D�s��1�듲��q��{x�����1�?�Wn��K�/8��h�G'$	:������j���qx>�M:���Ni9�E<�^�6�v[�qm,�\j@�}��À�t$+�%`3��
���l�(�����Q"�)��s��R׆�E�Z�S����],hA��k�w�� Q=�Al��%y<���)� �x	�/���)^�&�;���Wh'NX`=���n��"�*��*n���!�;�4.�ɖ!W�9���F��\�jnݺ�>��m��O����J�3��O���|)�k�y�0/,�4}�������m)�g���I�����f���A%=a|�����;^�S.��A6��em� j�y�$��_��U�^R�PN����n�#��k$g:Y�q�� =�Зk�n�4��])wM�����o� �<*��YV�*����l��/�����&�a�}s4���0���E��48�&��rI��/3R2�3�ŬT��f���@$x��-S����n�"Ϊ���y�RzFډ�_�����5QpcQ[Fhֶ��q��HP��1�����E���GC�A��(*٨���Z��_�u(	+�iqb �o$i؏�]|�z�7�ḠLs���.u�#����)��'!U�+��{ ��ޑ�Љt.��{��DU��
�-沁�(��$�J��d��WG��[��3���
Y���܁�#3w�|��DN(�俓k4�%�x`��\�@N���b ��EFc�z'��$�GK1b̵}�}Q�pƙ��o��n�q��X�~+��c��Y�3��kޘ��l+i(�w0e5���w���'l,� \(V���� 	V ��z���XT�4Ō�g�Ƶ�%��2�������i\���v^���'�$F�k�_af��c~d`�۫X^�����q�S����y�l�o��u��`V�ٝ}����ݛu���,3{�X�J��&2��_��g�"�Rc��أ����Xo6i�$[����Tc�\��{�YyW��0R�R To�gs�}?�ޢ�Ҋ��])n�6�8�h��Ci��還�3phyH�R|����L1A���s��@|u�d�iqc'�uٔ�^}��Y�h���sB?u�T=���&}�_6����_��1�Mp����MD��n58�x�s����2=׬� M�����t9�k��a�r��R��-���2��$/�_�rP��9߁�	�{�Q}#� ޓ1\י^ȓ��v과l�Z웕[)i�e�'��{�Q��B�+�K�߼��5�uKå�_Q8X~�>��T���~���jD�����?Vf�N��U�TC��]�?M���fge��	
���|݇�v\G\J�'̺=�:��>�Ty�ܒ�i�b��j�����(�qQ�ݥ����kE����z��@�J�.�e�S�2�U��f�t��F7"���:�0�h,�9�{�K��<��{�5���bۡ�!_�>=_�����EpP#T3p�biW
�(q�贋��#r/q�L�XЏ�鲐�,��㼾�S�6/��e����{�[�(H��*�e�D�;)��;K�G��?��a��jnq^h��1���i�k�b���-��w�4��fd����1+3�6%��]}(���5{`������qP-Z�O� X��YЫ��e~Nx%��E�M���RB���\�����LW���,�@8O�Eiv��O3���O#~� �m��3�*��־k=x��[H��������V�ض�aXӡ��k($>/���ZJ~�ۊ�1�7t��!��쁮$?�iJ��h6����`��:Aa��ELl��O��Ť��)c+h�=�龰���JV#K���tPN,å������b��PH�c8�_S��0��2���m���oQ��jޭ�q>��'���֞��.�@p�_n>����ls����<�o����
-�M��VD��\W�w�LV�o�Y�'P�t�3�d�<O���@|؟�	.�G_�� uIμh�B�ëҜjQ�Lp�	`̉�� K�(��g��_gg�G��-<t@��G�	���S��|V
,�LW+1ty�B�NY�>Y�$m���8tI&N�tA^�O���nZ�o��y��Q[���
2}��(%��i���z�c�A@UV�hSd�'��?p37�q�t$3e�ͩ҉@�*C���en��Jqp�t6�j���-ͭćUou��i4;] "%`�4��A��jMȓ��f��[�;_b�ϿeT=�w:��W#�8�1����{|���e�x��'B��v�����E����2�]WV�Y�]Y%���_���ݥk�U^���}�8��e��k|��<F���
q��֡U[�'})�Ն�7��}x윰4��k�g�;v�a�͂��A�yD$�uU�8��7�󎍬^`6z�'z�(�y����Ai��>�G�o΅CI�:�1S�mӏ=��0���nx�"�\�̕
0�^��������)<?��LJ'��v���k�mfK�-�H;��V1m�^�����HL_wq1�v�����%���(x���+��A�G���k��ydM�S�iD��]+u�F@D����ʂ��??�F��8՘���	 ���$�D�Ž�q�d%�qiȁɘ��OƦ�;�tVؾ�Y߁�*��N��53�����i�G��o�V�U�;�)���Z�.x�X�̅WX����s[��h��q`��M�6$l�x��V��U �(t�H�=��*��B�n�vU �!�_��F �|�+Q� %����=|�ٍ��m^�9&ƛG���>�����
D�#1�Э���x��H�V�d����]9la-H����ii�G͊׳�4e��1&
����9qV�V0tʩc��	�+ϔ�2�9xJb+^��?���T� Py	oۺk��/R^a8L�$R��ђx�l�)��^�A�?���\,��N�����U�?�{4�,�R�$��$��'�D�ȥmK��ndQvu�Ĺ��m��Ca��u@�������D���0�)ZR���K��^�n{��lƲ�'�;g��:��S�@I�Y�]�Y��[���aG.� :���$k`�t���Ǻ��/��Eyn�����&�l��*�?�����dzm�V����d��s�Z(��P�Lc~���`����:����	fz�0�y-��o^,��(