XlxV64EB    fa00    1ea0�Y����
wU4]�I�_�6qX`�fK���;�I��Rӛq�������Y�v6K�c����pŐ p >D�qx�P��nXmz�&�!��bs��>JM�z�3�3 )��|E�P4n�_��/���1�o�1�Ɩ2/j�@F�u˰���dA�ɋ�a͋��"�4���b�%-NN)ٰ�����2ḛ��}]�k>��/$�k�<�'���We�������vд���@�����T�(2��z���a��$��;r�]�b���	3�ɉ��*���z���%�0�HW�w&���h��P��:��$^�j�ϟ�����|'��m�O� ��	 $�^� b���o<&�14�nl�	��T1��K<��ZP��u\��*X��r����(�cZt�^��;��~�~(b�O�~+�v������Eǝ�I�����Knd�-�L���"�PM�����y���/�y��7�;�((tP�V��p;p�v_+������d~O��I �)�D�V
60s��a"l{��[Q����Y�H��G����q�F�l,H�0!�̤es�g=r��-��0��y�8� ��'�s���;,싑W���v���)�ȅ�H�
:��� �>��Jrj�W�vd���o�5�<m�� ?5���y�"��SV �T������e@�*I������4 �l�R�J�1~2�J
B����1�e��h%���Ǿ�*r>��q�=��m�Z.ɏ�����̝�g(xvb�v
�'��}I��Mc���ٷ5�Q� ���p�fq�V_d��=�ojA� 5t�#Cn���H���3;4w@T�V2i浲�� ��<���k��:�j𒥹� �&��n�a|ٛ��W�4X J�=^�4�=���(<�R�x벼�A�Ђ�g!={�)��+���Hø��+���B�D��7-�u����h�ȕ�~�wg��<:��ʘ"��D�~�s��u �#$"�o���S�����J���O?zW���\Zl��Q.�S�����Mi���|��17��L��%���;���^S��_q�1���:�>�
HW*�h��u�����-0���2��;����sx�b�P!r��D��p���#�H�.Ϸ2qy�J�{8{Àd�I<�x1�g��SRtɐZ�WO8���]i�lX�ϣ��~����
�dj����J��(	�i�h-s�+�"8���m�38xg}�ŗC5A�z��@�cb��4�c|�h�7��/b�Im�U;%h���J#���`�BpL˦ꤥ!�F�kֈS�yc-�K2��?_^��?y�'��Ng!p�oH"����g��F8�$1K��+��_�ݦp#Er�����HU��,徃6v�����J�w����Ka	%f;�s$��f����ى��+K���H�+*
̻�ߗ1���6��^�yJ�����_lv���z�{$�YF!d���D1_�����������]y����7�MoaD�>]QPsd�ܔ,���Ў7i	)TARq���`O5(���D'j�`�^���sY���5��j���j�E�n}<Q]��0��b���A�Re���?��w|.m�3z5/��X�{�}�i�qU��O9��n�%`�`�����Wq� :
�����U��ĜpBL����q���22�!����9.L�]��3����=��/�#�D��U:@��I����oQkڮf���7��u���B
B�����xv��rX��J�F��:����2�*Z-Eì��䙹�5�	Ld���v9��K�\�sm��kF�r}2��f�́�iC~��������J�u(7���P��{k�[�������)�9�{����]J��8zC�2
�H��]+����8��O�7΄9�7&r�4�UAs3ѻSzMF+��dy.�dX���������Z'75Dc�,�Û��En���n���)�ڢ0��Kp�?����!��Xr��C�,��
�r�2
bK"����]0�I��we��^�P�0E���?+"���89?��@v��^o֨�]oaC�ҹY�6ٹ�Z��Z��C�Ro�UM㙙Ve)��?=�JP�<��E:��t���G��,�%�� _��5�?����>�c��ۻ��H�&)��o_��ԇwڬ����L}����;,�1A��.L�e��A�LL��]<��d���~�8K�X�3z��h���r�W��9�eEU�Թ�ݼ-�x�!��"��M�\"���.�Y��9O�q�3ao�"��N��ŝ+fci�0
'���yu�y3�x����1�.Ћ���җ+�����/ê#��iYa�}��,�>�#��^H����.$Ufg�u��<�z�3�5������wh ���6�����B"4Ϣ�<=��U�Nq�J��>���X�y>Ep�e=�T�?l�Vz'�-F�m�!o�V^63�p� ��=��y�a� ��)�F|&����JH��6q�y�Ȧ��=����Oc�\������v�Y�ֳpHs������~t��)B�G�$Di�k9���L�����!5tX��t
�S�Q�N�9�=��`�
K�V�����A�T�G�(���7!d���N��G3vf����I}Ŗ���T*�/���n�F�߹3���>��o��u�FX��D�Q����;)��k����ݞ��G$�?��z�w�n��.β���F�J�C/��K�,��l�?x�U��ڣ�YՖ�����Ԗ�I���M@ϕ$�)��S����!4�ƪ
�<E�(�+:�6���6����}����Ɣ��2m���Ӥ>�z�&2�kM̦��tB��)�L�?3��� �����i���cZlo��0�|�y\�ȹV�fp�z2����*�r;��g�U4=�<�I-8���aZO@�f�̺���jM��?Ci�HZ��Z�A�GC��z[4�W�$pꨅ��N�7�΍�:�I	�q� O��:�oeB3)'�+��˚�mv4(-$6����ɭ���YF�����BwpQ�k}��7R �|�>-�a�*��*�8>��Dt�Q�Af�o��I���h��&�đ�;�rF�1�������&��8 8$��B3��e���`����8�7��T*�TC+zT"�%���BڌI-D������%^q��6Ƴ���(�k�U�7��(R*,�0�g�$W���.�F��6�8.���(�4�0Ʀ��}��Ds�ΰ�Ty���=�`i	���u$�FTJ{������-�\q��@;G�#doL=[|T�8pR�s@�LRz�޶����}N�^}"m��\Dim�wI9�~Ǐ ���D��W�k@�6N�$t�K,p<�8l�5�#%`I�~�w�a�/ES���e8���-���d�%�c1n	�]u��D��5�`�X��.	��8fs3n���d���g����+����vq��`�v^Qw�B��- g2t��w�P-�a��`���
�(�c�^�X\!����Vl`��zm�\Ǆ �2T�<�2N�S�LF�-��]ޚ� �� �~�����Z�_\w��6A{�w�:��=x�"a�[��{"h�� ��4Hn��PZN��Np���?�Y�#��W�ٰ�^��+`�����r	5�o!.n3�[gn��Ժ|倃�g+5�\�\�:=��].� v�p� ���ϪSe6���`��%�\u�^�L�Uu��Ƌ�w�>���2^��7@=ë�R�0����7���\��z4��g�KO0g#?��-�r��ӦN���9��w�@Us��a� t�Y�\"sd�>G��mMzJo���<~ -��_n-���Z��Tm`��R�<<iև�j �%���opO�#7�u��1���ӯ�۫GW�r�j���_F�:;�#�ZNzQe�PV����!��	�_*�}�S�ZxFhZ���N$�P2����( ���} -�Rub �&�݁��
�j��uK���,h��XKb0'�b�N�����*ç���}ro��4#�H(�u���6\������gv�	�w���ҩ�^HYs{��X �[9�޹����C�G�R��chzlUB*ks�S�����n�(����a�� SZ.�>���C�YӃ��� &]�P���D��2lliOz�p�/M|��_�-u�� �0��rR���Z�ϼ�+K��-�)6��2���8���V0{N�˜Ɇ��I��s�N<ɜR	� �Y�gQ}��y:�P�{�}l�Y�'呁o ��*�.�@V(��/�S˰����|�Vbݘ,_�wԇ>5Ž~�<1�aC.s�B�1�Ļ�.�NO��jf��L(eo��n��e����)�����ٝ�ksg�ʢ��?y�����Y
�n���+�����hP��Nw��ەC�۪f-��+0ܿ��ɷvJ���~��3i���y��[-^�6�\��9���ʜ
)�]�<< ���XAQ��ʲ��8V�C��x	��dm�0�hDt��+l�Z����B�L����x������l\]�#��A�@b���y��?��A���w�����9`uv�Ž�/�i�Q��zE8;-OU����E�lT�ɝ����?�W��/��A�,(No��8�d��I���o�����B�*E%V�|���~jY����e9��lL�D�C4m_qL����FU$�d+��.%_
򐃌V��;f��4�{�N��E�dΨ�)����M�f�g�.��̑�~�z��<&���9� ���+ͅA��Z�J-rl{
eGNwT#�����[�QFHL�S�r��1�w����8�ɞ6�D����x)�_T)��Yr_���L㤃)'���DE�.�b�)jJ�w��8�K��n�zL��"��$pa��W)ug����ƍ����M�T�;}�Ʋ�a�x�� �L�kAv(b]z���h�߃W����(�q ֚l2'a-��:M=aJ��P�U4�ܩP#o�5��f��q��ɉ�\��	P��P�g;0�����z�'�;"���A
Y1լM�pr�wK��ڥ����aV�*RO[h��ZF�D�6{p	�!��X)��B�(GSc����O(&D����Rc-2*q���;5>.S����g��;.Q�W2��C���{Ƙ>OV�#p�~�����9�P�0�_�F��[뼐N��b+.�_$uh�nǇ9�O��d=��� �Foaae�� P��R���k5P����&l<�)��:Ut~��<�H�|��p�6��bD{�aNG�'��+�<�
�Q֤�H����}�&y�l|Oݶ�u���+@��@@D�+���?8UI�v�^��o|�mp� �;�3)
o�_�-��;1��3���w�����|�W���MُÖ�����_Brv���"ۛ�4��ԁ��bsLMB!�E��Z��e�$1-
�z5e09~�oU��2�g��财�Aq.;��h8�d>L+D^��:4Z��㨟<B0n�H'&!�1҃4����d2�|�ԥ��p�;z����{����Ky,�������1=��cG��Ӎ�h4o���ұx��$���O� s+���<�/L��4���u�A`���=9p6_��SRQ�-�6�A�ke���\9m	Q+���7��Z�����^��%�u��P�L���W�Tl���������''��&�bC��!zH���b>J��i��'�i��{^�2��
���-PN��DyD��@�0gRm�U�z����N$)����Z�����r�١� ���訙����>1*U��d���2����!3�)~�{���H�np�:����'�j���z3��aT�$hZ����QǊ/�zj���Pd[+�X���z�����C�h�K�鉴�����6�|�ۗ�6 �Bu������ߐsLbC��f��Ǒ�D?�z�c�������Jt��א��8f1��|QԄ�,|�I��'ķ\��� ���h�i	��ʧ�f��彞i�3>dJ�M�$���5�trC C��o�� �1��z���(��%�'�b�U�.�6q\j����U�$�.:��[ͭ�?����*\�P`\4m�Z�'�{��o�|��?g���6uR�8����0T��|]�Lݗ�X��x0�S�Zk�b�I!��<f��3w�d�u{ޣ��0ۖ���T.p�4NJ��V�J�֍"���:�Uqxe�|�Hq�r\�ԋ0���n�\���f%������&B�L��[�LSٜOO7�S�H%��|������W�A�ޫ��+#1G��k	��&���'�R�t�ے���,��溷4��qљ��ڬ����Z8�H�՜�=uܖ�z�]�WIm�G��'P��߰�SL��Ȋ>O���Mb#�d�􁜤"�n-oI��o��WTRqOjۭx�'���I�/k�IQ�L�N��^�AH�Ͻ��aCQ�7��i��EO+v@*��.� Ir�����a"4=`.пt6p���ÄP�gkG��
_g�䏉[!P	8��ב��>lQ礶x]9{�d�SoQ9�t+_[�4Rx�F4���I�g�%��� =<���6�d?aDc����{�
eJ�"�ˮ?�<,B�?ʞW� V��P)�`���k��f18��dcJF:� �dR�6�f?m�v���4J���!��J�]2��=♞$�V�feW���Q1KF���}��ɯ 4�:�YNB��?̽��c@%����̄�d4&w���&wF��Y��=q��D���st��f����%�t�G�z��xo�"��l,��I�U�u�:ޒ��r�3���B�Tƚ���˷���j��&N���+2���"�CNJ��cpX<Y�5,
�����a��q�8��؜d�Y�����3�҃�%�kQ���Y�����7&R�1�|ů��^}r_hW�>��m���n��K�h�S0ez���%��<(�>dt��A��r���b���(Ɗ�h�+'-�����R��e=}�
�����aB7kW@��������;�ZwX�; ��B���*�Y� �8e�t����il1�}"̚����:&S��So�nt��V�B+a��'>��t}��uM���Q�/F�'�6Ri`����X�P'�.b/ņX���st����(+��a�E��}�d�Jj^�E]#�,:� ��)�ۆ����=h]!0��Hr1-cgX��$�����K:�Ɵ�ܘ%�L��z匕���i����쓍�<EɁS�u�;�A���v`���A�O�jP�plU�NO]�G��fd�gѰ�l�[�=����M����{;���^,�js2�yH�hp�Ʊ��E4Bw�_pn��&���R��8����f�6Ո��DA���0�
_#���m�P6��u���������6�>4.K/j�Ɗ[2"t޻�Ze��ГĈ��H���-[�}�~P��.�U5H$Ts�ݪ�ʽw�g�Wv����tEĀ�>��&iB���" ��Q�1��_���<,��N��!�Q|ꋫ,8N��<1���4xe8߲��I��b�8�Tc��o0���n��6��I��K\?Q@9�o� ��g�n͚>�P����Xa+K�]��2eq�f�!m����0�1���fB#O�8���G@���K�s3��^�BۙΔ ��b�WW�	��[sjd8)�`�B��c!|��e���l]���[�.kƍy�� �aµ�u���x�Uf&b��A�x4L��?�n1�.�"<�Ԓ�D�{8XlxV64EB    7b11     cd0�:��VT�+星���"�K�P�������4a�������W��Hj�6�4Z�DЕQ��jVz6��"V�
b|��u��EX;�".x�P)ߣ:s�X��|���h���>"p�	ra��~��t����E���^��JU�\�(�g��hƿp�X�O��>	h�{������O�~Cp��/g��fHXB��|� ���#o

�xWL�j���\����ڊm7niL��n��$5�X8�Z/�s`�]^Νg>;6��s���.�a1ьtS�t��	u��g�f4���`X�  ɮ�5��~`O����,~T�������GZf�\� ��<o�*i��� �B����y�T�DU��FS�5�6\�ۜ������J�����P����
��F�*��T�0n��p��I��ek}_d�����```�x��iP�\m8�)�[�֛����6�E��<n,��iއ�w"�M(�ED��dȹR�������E.ɉ:A��#�u�+^3�'%� ���_�C�q[/��/�P�h=��Ʊ�!�>�@D���lK��T-�5!e֖7bŰ�P'�e4�A0&kܯGe�s)ǰa����ٝ���*�l���rTP��\�4:6M�e�R�����Lh�>�Ubĩ#"�+I����Y��e-�a))�� ���$r���0�;�*���\�X�k�ꭴ��y'ftk���@ �Vtk�!0��ޅ���K����n+��P��*:�[$V�R��Kż�z}����X�Еi��B.��)v�D�E��7A�_���[�/�R�4����*C��`͗�6C�����\5�yLJo5�mv�H�� �4H��
�Fqu-<��]��O��GyԲ2!'�f�*o�5(��N�vTZ��Ug�ٶNP����zJ�� �Q�oD���GS���&��K�tZ��U:�4c����i�[َ�1���=Z���|\!�^��������]�-wȩ�ā��G��/ �6 �X���=�ƺY�L�$H���F�&��Uf�C{,���.B���T���Z Щ(q��r�
.��;�=��=��C� 
G� 
>�t��g�H���+&������x�؉�#���^I����"�䈁Q�	�p �팆�rE���'z���F�����̝���<�z��>a�VDim9�CK��鑦@Q���e��l�A��[VcBd�'^�E^��o�Cc���t�I���Yp3�,��K�k᪞&�����Hh��~����h���/۹�`P/
,�(+t���㡑z��K��^g�,�D[J�d�������,��r�^5������<��q��h�����A�\��=���c]x	f�e���5h)���(ԁ-��NNԤ�Hy���|9S<�Z��C	*p�h�Rg�U����lJ93�T��7o���T���/���5�R�%:���z=�	�e�j��VxN���>���$bM�2^���i���_�3t#��,�y��y�e|����WUg"�oS��8:{">�g����vh�ᆲ�ޛ���`͌2~|L	�޳�X�MHxJ
��gB�}�-IeR\QD���mj�i��#�����c�u�x�#��2��?xH��u���38e6�uF�2�3��I�!��\^j+��.��C�&�����m�۲;�������%�^������Du�ǝ�mu$MK�˓O�)T��t����B�ү��;�����L��{�!���X���d���}�o��3+���8�0�q�T^H��~���SH@�e���Y�ݹ�YZ�S�������?�`Z���/,I%H��3?Yƫ�xmC��m���(�;��>2���`�$�قM��oN~�6���<���㪽�r_�\�6����3+^��;F����2�\Cw�M� �����#�l.3O��nX��v6aG��v2�`� G)0%���q9���*�c�e*)��,�]��-�����-\�-���^r�Z{̔�aU�8��4��NB�yzfJ<d�3,M�7�g�@���AG/Y�$�7����EK��|@�T?�^�7=��
 tK H��^�E�,AD*`/sQW�d<������d�m5��yy��S6JC���Fz�R��ѯ��tf���I��6~j�X����p.�m�%��!-���3�ӱӓ%aS��6续���2zڬ�H/�����^\���}��ؗ����ƛ����yV�F�d �eGϯè���oFX���Ԣ�
}��3��ѦN�^������!�ƈ�;5��TL�.J�H2�e�Va�&*.E	��5�7SC�s����%�
�&�}�����Yo�.ʀ�Q}t鈼ǝ�b�a>E!(�{��e�ކ؇l��i b`��Β�a��d�Z��;S���H���t�[��Az"���L.v:�1���y"��	��R�(�@G�&�����۬y�)�ޅ'�����TA�<kߐ5������Z���s_4��m}��g�6����G�'����,?mi�^_\��٠��r�^`��_8��k3�}��١�ͧfg���6Y���5�)��K�2�;mGE-G�J�����p)�2s�ݟ`���߲���2�"Kr���w��NӴ�ɛ�0s���� ��CH޽u`�p���7�/ؼ1d�0��S�W���s,���=lfǊ3O�%/��Z@Ƥo���e�7��K͗�a�a�;n��H6  �g	4��T������]�k�;ۦ�B}&��s�/���{��s��m�*`���}��=W%7��/e�j�����m�~r���؃���-n{��㦁�
Ԓ�ʇUTi��׎OٌɈ#�I�����p��a���L��̴`:%���0���ub��g_ћ-� M��z[���I�OT,�_&N���*���q��?dO�o���(�"!}(&t�ќ������{��3��0�������;�:����*H��(���KL.��O�<0�L񛄶䲰V��
��0�k�(�̭wƃk�)��%n����\E[�	�nZ#iNz2�O�٫K*^s�RNV��+���%���6Cx��\�'д�ΐ(�H�^M} 9�(f�<�����ߧS�"S��)����L	mפ|�X��r�_8u����R�wB*4��?`�) �*��ջ�8��M��>lz��E^ր�AS%����n`�� ���!�ԯvJ������$r���&A��9�l����t���d1��.�0�;�5o���