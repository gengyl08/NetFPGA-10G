XlxV64EB    39cd     f10.�k6	���wJ �����bw��
�7'�#�&۶��I���VM��&��C�]�C���*����>��h\��E� #����qM�)'�u3��.�5Y�����-�Q�`�}�q_�Z�d�����Dm]f흈�h�ټH��vg�c�~/�o�!�VǅV��%���-����ž\���r�
+lA��*=�lB�+Շ>a��'�)4U�do��{����j�Y�q�IM���j�˛?c-�>���i��ծOq�����^:M2i��M؉�m)����
�dI����$�_�4M�v���<�������@�J9�bh��$v�'���l�d'!i��;;��c����NUnk�����#����j*��5E�R�G����柮E��i��J�+�ת��e]�D��}��j]�~��X>Mέed��D�TK�R�w��Z±1et.��|#����׉2����_��.�	r�%�Wo���/�SФLÊg��0� ��[ID C���/4t%�灡9('�7��˜V��t��
�g4�OK��ômUp���7	<�h��� g#Vj�2�Ȗ!��n(��bc_�n{���'����n��c	��4�'��r��]�r�!͌o�}�OB�[�E�?B�k`�,�]R��d�Z��]Z�+`I�?�j9�12���� ☩�$B��hgڮ<���B�������
ÄD�4�wseu����q2�@4ێ�`>6����"-%	GMa�2��}q�*I)����E�%�8��d*<'?�sd���G��0
��G-q$Ō*�#��uA -�Lt���d�q�oO���([I`r*Ui߼`�?��3��Lz�=ݔ;Ux̋�#6���_�A�^w��u��esC�$��}X]y�Pݍ�J���%H�/��Է�*�_�I�>��-����R���_2/DN
�<%TRw'�:���D���!�B\��}ˑ=t3�?vL��<W�Ym��%��aC����^�t��n�G{�������6?Ԯ9����/3��B�����x=�k��3�O�(�ꃻH��9���I��[��g@��w+e`���P&�b�Ff�k��=���2�pb�!�� ��c�n�ܲ�w-��B��U}��=V�bF#^�ϣ���X?D�<��ú�\���=�<���Z�%9��ϊ�9 �'8=����L��@q�m`�T�t��=��{�C��rm�&h��D�g��LH�B�G�������x̤)�Nn��:�=W�l���EcY'�ܛ�.�Gک4 �s(�I�E�Ҙz��? �\6�t���EM�ܞ��m�F�zQ�>��|á�_*�a��ы�!
�X�W@���i��h�����X'|/�[��G6*]P�(��h~bu�e<94���ɹ3n�y8���R8�-����9�d��]w��9������+��@ y�Z�|G>ČT;2O
��RR�j*z��$��C�E!/�O4��l��I���1;�U�Vp���AE�TԔ�z�ޱ��L٧�R1#�W��(��K��Q�9���m �wx0=��t�V�~�� +�Q��N�\e��#L�y����H�t>���/_�Z8^gO����7:Ϡ�bq������i��NgF�8��"��ٖ~�}wXA�X����G������<G������O'��Z���'��d�8��֥UfN�ΐ9�u��;���y��3d�!?�h`zt\�Eh�T���̰�0ki$���p	4i|%b��'+^?���8�k�a�Y>�W�ƺD���4�C,��v�'�v�Q��bT$�}%�rfߕ��n�ڠ�\��R�}[��ݨ���T��=]w@&�
�$�_:�}�Р�(�����>�-7��&�}�f�q�l��9�Wg�Ւ
� ��Έ��� >�&��5��2�3e������}g�JZ�
�S�
��R��-���Gr����%:g]�L�=Ћ���?
.�`����v��a���P!�h�{d�l�ن\3� ��F���-)H:ɠ���U{- (�f���΂�Y�Z����?r�>�R�8)�2�j�ˠ���EU��l�tQ����4���h+� �k����꜒�"�'�� ���P��'D�Ν:ڛ��}k�����U��.ǑO��L�q8��'����.'�xfʈ�a.�<~l�]gzu�,?�c���`x?�yXBr��lp���L�8�f\�ΎiB��^�4�`�^P�Z�C-���Z�P5�4tCk�!I��HēU�5X}���l�r�����Qp�EpAs��/� E��������Wjżr�75���Li�_���1	"��M�6������ Tc�.�tZQj��d{ C��1����|�p�W!��Yv�` �w0�muO�@��n^S)4�,:�e�XW�pd���c�WO�HE������5�?�Nq�~@�م�@�:���}[�o�Tꑏ�;i�)�\$=c�%�D������@��<���������
:IͲ��@��I=��WQ� y�=/L?�N��`N�ف�D�|�\�z����]8���Q�!e��E(��B�����Q
gC�p�����)�2ޘA�+�C��vp^�8�[�Ǒ�$v����!����7]b/��j%^�p>#!�~6�n�߲NۻD֚����ᆞ��W�i�G��i���s�~�L*�m�\*7�Dy�R�����NK��:��"^����	���i�ԥh�!�I	�T���_���mz4[���fa��8��nu<������i��`�����V:�,I��������շ��?�B'{:0�o���f�,@J!�3g��
�����٦�.��4���g?`�S��w�+]�Y����ZU*)_����jK�t���A�Yr�.�`��6vAq�!Tڝ!���T����B�Jo���y3^M/)���ܯ&�d�XH\b7(���B�!��ƋU��1��#��jɗH֬kd<ʊV�4��96��^%x��Mt�5��b�L�.��)�s`���Io>�e�'\�~V0�u�:�#>em<�6��j���i���M]À����L��5<&!���
�����U�1N6��/×9�xa3���QW�>vg�4�a��i��������9R�i�����6�Wi"+�g�g�F���FP����P�PY��S��_qt�9$���4�Q�o|_�����;��WXe��>��dd���T8�U��^Q��8�ڄ�Te��\je)Xy�jCr]蒈��r)��zTIQ�[5�ۋ�!�ʭb�;��	�8��Ƈ��j�/`�����M���$�;����V�e��(��X�>hXUQ��_�	�@���ML�SR�]ֿݛ�x�R����G���X�ɍ�jN����]f �Ǯ���U�d�����@�y�*رh)Jc�~G��~0��	mj��AT4��#Rb��rX��4�p�p,[�D�h˛�ۆK$:��2yr	)B�΢S�/q&��l��hv�¶�9��9.��v}�t��d�ƥ�5���1���w ���y`�tkC;��#i�~�z�6�Ҩ�&U)�ˤ:}��`>9{y:e��VM}|�T��.-�Q��+qF�قf,gc�cc��$)�Ű��0�o�p�g�:�6\j(@r�z����Ậ|���V3J�w'�ޭC�,"�s��9�ں��"�h'GlI[�;Y�M\Eg��&T%©��J�.��˓N�'�Ʋ,ag�?j/v C�'ga�8������b�Fv��]�����Q��|���CB3lC��S�i