XlxV64EB    28be     be0���4�A�� � �qY�k-"2�w[�&�2D��?�ϙ��v���q���{��w��iR���� \�O�2.ʷ�D����s�Bf�^1�OS�7}���6�m�� Qv�z��<��ߒ��3(
]sb�FH�M�3��V��ɯ��ש�i$�)��N)\�T
��ķ@���e���H��z��(;���x��Qtߢ�,kC���A�M ����a������&~=r�$�$<͌�te���k}^�3i�{5�qf>  T�c�'\��ZLz0�_�!q�F�Lz{fڛ�J�W���gvU-�l>]E����$5*�q�J�*�B�r�!~����v�0g�M��mA#z���7�5���Qq��2>�?xI��.d�&ޚ�8�O2NFM�S�b��qH�`�،V
�|�q~[!�I~�%�a���j��w��I���u%���o��^Ջ�v�*��5�w�M橛; \�V�Ƅ���Χ��Lh��r�Ή	=�z�*�hx�,��#wh�UzCU)�Ptˉ�ey�,�aM{�[�%��NX p�ʜ[����<�z9����z��Ci�n�P�w]òGF�����H�yոY=~��LٵwÇ-�]\���;��0D8�:Z���p/��:QX.����^��nB���tu^����c��x�1�		�ý�eR�P�����T�!5@���� g���3\���>d�0x�0�:��/!�<%�	o����sK3}��\���}�ƪ{J�Y/�����!�D�ce��zo�x;�p2.+M*jSN��0\^�1)��b�C��T1�I)�����~��T�l�����2<0"SܐHK+ynf�jC�*�T����[Cɟ5�D���2��{��|�����r������'	S��M�N��Ozb�>y��0���ބVw�T��nւN����ok5�q�.�Oq�	����z�(��c�[�NvS��/%�=+�ţ�mG0�@��[0��y&�u��_ٴ�_����{�cR��W�������ȲwhS���HJ�Q��gy�b��� iQ�X>��:l4���/����:���+��EVka�<-�����ǵ
էt�UN*JK3/k��}��E�����V~O��tO�k*��y��
�ʰ�u [ӥ1r���셺�->N�Ȅ@.��0��ik�U�]�o=��d�0��Z]x[#��#�-,c�l!�ɢ��+c���t3�J�Ha"Q�}���A���A6�L4e$�ߖ�=]-���ҫVc�Y� {`s6�����+��zn���;�'2����g�Q���|c.�O��):�D�|ԫ�$-��\�C$���F���	<��F���>��#U��Jj��~
��T�8���X ��1nf�u�g��uߋ���$?���N�*Ԅ��xA �W��%MX_��G�&}�����R�D�g�"R�k�c~
gN���9�$Q�Y4����`�o�ۛ�rY���*�C�B,���0.!R= G;��n>�zP;�1�GU�	��Ç@戹�b�V�����l�y��<a���i�©�Bx�����j><�L�I������2݃/��{�F� ,��3 R�mA�?��:,����-�:Ip�L�t��:�9j���3+�� ��s*t�+'/�/�B�쥤��܉��P����&�i��j�Z��O-�G�WNx(5*�T٢\;�B�G����,*����ůn3���5�/y�.�i|�wۊ�Jᄭ�Bh�)�w�˶�
!)��!<\�5õC��cs��.Z�]2����	Zp;�ﱜ@�f��
"#M8�o������N�ޮT���4�H�$3�#�.�h�S&[ٵ6"�MN�M�z=���ЎS|����s`�]T�$s_���xg�oa�XC�Խ%sb���:<��Ѿk)����.�'Fg��/�F*N;T�Ȫ@s��p��l�,����n�@#��UJ�H�����lo���O��)����*��W�5�(IKP�%�%Y���%�
��>ɵ����15/�}�X]:��DaПL��=���,�K��(e��.��B\)	���/q������j����/Et�8��m��D��%4�:�D�Xה�� ��v%��T���%�@��2ͦ:�'�5*ճ�8��`Y����CV�v���<�/�/��=��ީm��F;L��J+�ІP) y?�����7o
3Ιx������B��p�a� 
o�9��3��0~Vc5&�]Rr׿�$���kk�,]����,އ�Im�����4R����=ʽO?�,��#'�Loɥ�:�Gty��:gC�t��˶U������FH�X�# a��O�]O7�W{�+`6n'��h0�9�1��[�5�Ý���*�\���@F�
�p9�����j��_���i|�[<=��ϹYQ��A��E��:���#�kE'"��.�A_B�8-�ԉ���k�h�۝J9u��5Q�U=q�Bdȯ�	�#�ɦ(CyP�鏥�K*de��ő��25f��De�ۮ^¹Ui/�!ҝ?P�j�&���>s�����7������C�P~r��;Y���פp���I�ag$}9_�4�EM�R�͗j�jt��Qeq#1�/ɗܐq�y��|@^cS�%.}sٶM3�B1�ϑIɂ��1��&�3]���/ g�U�ZJG�>���.��u��2��Z�E�83?�1�h�gk��إ� >~*5¸�L]fL�]�{��2-�B�g�!��O�{n�t�u���cF:`�Ňt��b����ݥJMGwǢ��_%s(��&�t/�� a�O\��E��+�Sg��mb�@V2H������k_W�b.m��Q9���>sx�.�����LzZ���A`el 3���SѲ&�m��{��)А�R����n/�Wт��Ap�3�G9Hz�Y��������#��wC�압��	���OTd8�üֲ"?����l