XlxV64EB    2a70     cf0<`�0[�����i�=?�a���Y�/O(�qR���-iQuZʴ��,(�ow�'�t�[�U��` %��u�J�f�P�BN�;,���>���lMc�2��t��U�D`e�ͯ�bՖ��b�&�ߕ0��2mT�=2�`Ճ���L\!�lZ7Q����%�wv�:VOA��6("�RU�Be���b��\��!'��<�o/��f��~�-!��|w1x���,�/q�z-�kс�%���H��O/�/g*ƾ������zm,�d�ď�e�����py����[y�P��y-��Fz�T=a�C�%f�k�<}�O,�g�| �t�.���*�G�lv��ѥ��98PR�z؝�K��י4�W��Z�?��mo�K�:�וg�y�
��5�A���0�Ο��6�w�g��Ug��T�e�+�[ZEJ�@��m}�g��HW'��Q�F��O��͎~�O�6=n2�#�}	�}l�?��Y0�c��*�Lk���O���!X�9��z~'����g�#X�����eFZ�A.!�ۼ�H4�觋fȃ��㪸V��j#IZ�`���R��e` ��DP69Nlߎ�qOȠyw"��'�9-u�{�"��L�3mcF̸;hr�n?f�A�l�;�?fLX;_h@<�zc=�a6�O*���ߺ��?�)�8S~�kO���{���D���'��i^��i$��4��Oy��p�R�����o]�2D s�]7���Z�"T�]�)�16{{�̎:D�ۖ8D�W��:�w��.�YL9d�U�Iۿ��:ܣ���/;����\6��Ű�H���Qh��/����xr��-ߒOሤ%��P	���ч���\������sc�lʢ�K�,-v��d.�9ȓ�hEٚD��k��:*���o4�z{��i�4ѭ��ćA�q-yC*ww�s����<9S%���D�?P9�`�P����ƨm�+�Y�����ZT�?`V@��ڭ3�T^σ*��Λ������ �aHV����L-ʔ� 	Z��+�̷iO�^̠�ǆ�zs+��,,����^CK��X�޳5P�I^���M��B,%�e�)˸oc�^��kI)��Jef!�2��r�I\�	 �	���[z��j8����c�RÜk�!��=�O������x����� d�@ ���c��g�I�Kx��+��$69EM"f��Y|���F����&9DJ��y�O�S����7f�F��Cpa��(ܽ&�����'D`>�G2�#l@�dNVs����5q��o�M�-]�W�<'��+�w�W\- ܨL2lgG�@rӟ��HƇ|PCsJ:/0�̢�G\��u��`vQL/2�na��GP��}a�ن�D$�J���z��>�����r>�x��J�-���hi<d�U���=1���w��|O�2GЅ*�oSR��>W��Ű���1��JJH��ZZ��1v���+��-�Y���l��S�&��:�~�czc`�ܒBe�@Ju��`�:���#>�sd�"�y=�e�p��֢�X�K��Ő�Vg��.��A�����@���P�ɕ/�a�Oz�&��ܼ0���p��"=���=��^�C��}����4I��*��R�Bq�<,Z ���[�[���@H���M�V�	Q�b3���Q�Ҹ��
�O�^yi���q��2,)��0��n!����R�B�����^�����T�T�TN���w�p����Ҝu��.��t��V�v��r*��Dov�F�dNJw�k3�풄�������pA��#@���#�T�kWX@�a���d�[���y#�<�� �,��;(i���ïȪK���C�#�z�ɸD7fV�8�������� �S����}�f��ߦ�V��vL����X�k��ѻ�g�j��d���T�.w!����rc��_��B�Ώ����W�2��o?�3�X��E�}U��]&赀���!�R(�IJX��Z� �)^�M>�yM�}}\��v溇�t��R,���7�Lʁ���'��Uu(>|�ôz(:��,�H���X��^>�v<�l�+��D�S���NSZ�[7XнiKf���0��)�8{ǯ�8����}X��`�lЬ���0��慊�����@�%�*%�	�u� Z�m��������)�X���)))ϱ�̉f m�S��^����B^���Djb�1��Q���͕G�r�q���r�NLM���*7&��s3����դ�V�\y����}�i�<�qomʇ�bj)��%$L�z9���_!9@��P�o�K��5\@ώ�D?UU�G
�!�������ĵ=u�� ���W��w=�f��U+����)�!T�9l���#G�]j�'vǍ8C�F�����ˆ^�z�QHbrJ��{锋��c��LS��)f=^�0���$2U�(��u9E�m��z�u� X��<�>	�����&u�0[��$�"�J��!?�c~3xg�W[d�{ؗp+V�;�h�mr�.i�,�p�ܷ�i��9Y�nL�[A�d�5Ŵ=��b��$���Y1��b���o�J��2<�{8�+�7�#H4�!��5�LW�8�|�Jv[�0���\Eʐ	����)����Ԛ�Ro���F`�,PD`O�H���[����j����9�[����k(���u,��65@��`Q�7|�-h��7�,���N
�q�eZ3�E�˔�օ&ַj>@��β�Ț*4�Y���EJ�v5���k4g�>����riP�)��#��]�V`�R�[��_iY�]��}RW'��$"���F�
��k���B}����z;��g������W���8���EY��4�x\��#\��Ŭ�)�|7� �y|j�[�6DY���,1�ԇ\|�q@{RRi�+���̺�n�	݌/Fn2�2nLd��S�f]����T�0�v�K�2���	��v�!�t�iޛ��f�g�� ��.�a�d�_7��P�Q%Ŷ��q��腪��\��P]{}�-�k����������CcBS�To��ѹ�G��c�����E�l�3-���-X��[x>Oڹ��Kw⹨H�B����'�?��4�:}C���,�*�j+�܈ңf776�����Hі���L԰ 3�!U�3��V�>�
�K$s��a��TSP
b*�]�͸���,���4�S_�{�J���P;�kQ4Y��_r-ݽ3�F<m`4��X�!{��m3�%��h�VJ�¢�7F&ǒ���B7WR4L\�>I�|�S8���Ӕ���N��