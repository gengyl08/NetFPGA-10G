XlxV64EB    b8a8    2370�=V3�L���,è����,k���J%��K(��o9¦�	;a�'��z�<O�Ku���1aӏ��D������cx9��!V[V�2�d�2�l�X�NF�F|�Y�N6G����ۋ�)���-H_E)¨�E�H'C�"k�:$b�B�Z�=k>��W>ɐJaWfi��D>Q�J�%o�/��#�xF���{x�AEn�C�m�=�%��|1��L��~�?y��J�D�a?$������x�d��A8�����>�}x�d�L�q����N��Y��W5Fs~�q�;>1�YLŋ7ɻ��r���*L.�V	�a�)�A��4�D�Pr��ҫPv�������Ɔo�C�pcs������q�G�������~ľtw��-L<�&�[8�Ӡ�:[z���zk{��l
��=;q�\�(��&эb֑�ʯ{��%OҖ.��ū���m�sO�����N&
N������/�B��P�����fT��p��]��,8��}�*'a)>��*l?E�w��)'QΧ᤬7���C�����〙i~�1F��Jv���m ҳ�&	w���_D�;_�U�:�@����YcWp��g0?o�-��V��c�W��[���,V��ѻ���N
?�~�b�)�t-FKqȽ���}�\��0J��}�����&jv�"|�R�MHƾ�3�B_'ľ�?F�ˠ-�
ԛ�;ӓ�����=�S��`C+�.��B���@�˝�Vu��w
�|*1ܰ>��q��Q ���n@��~a�����x�:ϕэ��b�|�K#8�[}q�g�!��L*�9��b��L��R����c���o�c��cpD�Y�+z����\�������.���2�$ ��2>��`��F`P9d����AHQv�%�ЁNb&���\mj����-��hX�v����9�#1�tV���t�͌�r����}S��2��y"Y64~7��K("�9����!���cA�Z��3M�Ѫ�[�����"H�ë*�B�A��$`���90e'x�67��+iT5�8�A
q�z��?C����M��w�DI� �$7��hW,����z�2(�_���/N�r�/�K�K��vj�q��p �K彄���=_Z��0И͂������"j�;M;xo �?3bY:;�H���C2��?6���\��cIk����P��b�Җ��E��6�><$HA&H�F�I�=,�W��|��F��HExh�P�5�z�w�BȾM1�=o˱��*en*�+<�z���5på)��� � �E!Dc$5ԋ��kf]l�Z��!�X$�b����de��=fr�g�#Q0�^ߺ�@�.�ҹK��~�Gg�~Yy6-�R�`U�'�c�,.	��Z�4�?���P��o[���1�0��8��K�O�r����0���4q�H\�a��I�TkR�x&�7;^>-�;�q0��(4[�<��Ƈ�dщ�}�vE�ܵ�_��v�PKx���q�1�������
ũz�ªp��ϼd�B#�lh�&_��^!�^�Rk����T�`0}e�W�r��gV����a�DM>����v0��� �H�i�Ӷ;�W��Cl��３��]6�I��v�Oaj塳f��#�D��8(H8���C�}�Ac$4�Ngz����9�,",�T1��n�t{@?zd�RKY#�@�.T��R�.�&�K���C(y�W`��,O��ό�7<Q��\ƈ��K���������K�6�^怊	���	,'kJ�f��	���������H!jD��{�6j�N
~��Kŷ�?s����n��)��6���?��iQ�3$�M��Y���?�N��f"�X͏Kw��b�T�h�!�]9��k��%,S��D��Tb�� �<J�q"B�t6f��B|^o(,�D��)��Z<��O�{?䊩;J����+ �]Cn� ��n��73��̊}�uQ�lk��MЫ�M-W�Tesi��C�ض$�n6��t|��3`���^��u!�m��|dX�Γ����C�̘u3/ݿ,T��j�\�����=�Ȱm�9C��VM[�il����
F�#�h}_�r��(b�p^�:�B�������}L@�M�\(,N�,�Q�-Ō�ƅ%�,��z����-�Ie�G 0���Q���X��i�,B1�9����e-�>y��Ǫ��z*�cp:��Fp���W��2�W9�E&����p�3��ヌ�OX9&��@L��K:���) @g��Ã;�&�Х�6tN|6w��0�D��![GbFwE���fCc��b�gnFX�{����%u��BCIv��p:�up�I����0~���lU_��y�N��۪lZ�_�T#�S�����Ƒ ս�����?���}=|��̫���%q��j�PR�<�:�p�A�F��u� �ze�ڧu<&�!v�IU���s����o$��P���.O+ɆNgH���1�v&CxQ]�~\d�\�Ќ'�
��_�y���|�O���8id�t15�X��CgFʹ?znow{���X�	Q�Ʀj;�M���%���M��۸�R�e�\7v2�K��4~�M:��vz��w�T�5�w�=z�����xlإY�E��o](q�������6��\�%��I8��Y�Mg��f������>Ϝ����kG�
�۰�!�c�Ad0��,S%�� �0��*�cJM�(��Ń������U�;�d�
M���3IA��v��^"� -�AG���|QD`ů9�~�t��pI �C�� y��-��}��(3��D �`�=��ᤙ��s�;B`�W��݋i&����*�=�G� ��j�.����<�?y�&�GYϠz	�lã�m-�<d�!�M96P,�JYa�UFJ_}-&��e��gZs��E��ߢ ͠o_�o�ά@ָ�	�W9wn�i,_�!'�M�Q�H7��E�6J�ё�����͸���^e��B��؆��6�%���S	M���~�b�|K#�E���J�?�E�Z|B7�4�X�d������2������j6~'^H�nC�(P���TzG�L�.?�%.h��xǘ����͙��0Yt�F'9����r�?��<H��g��1�7x¸$F�vQVu�W�eg���8B�|=6G�3��P�� 0��C3�뱧��*`���/>Izb��s�&��/����r�19��A����j�g��B��ٕ9x�#���<u�e�~A��J�p��
�+�$H`u����T�>��`��Ĺa^]�X�ԕ���Q��o8dB�%k}`�p�NKn�)-�$vgmh����M�<�p�I��剾WSܭ��ҷ̂,�ׂ�.q�	�;�Q[_x�zB�$�aKpE�
�ܥ�_q�a���Л����8O���r\�3sE�����x�m���4 ���V6e3�Y��IW�FZ��U�{�	bHn��V��m!B*5HGlB�����O��ת��KC�f���9�Ma�	�U��?�4�#���V�j��XN���S9k%o��&.R���?�1荷����l�6<�
��XVY`rN�S3Y0n*�z���o���~��bԀ.}���03�27I� �l�e>|�Hy_(/�D2Aot��y6�9�j�i(�$Ҭ4��l|Z����=��^'���mP�10?�&u��|`��ð*e
9K8����
i��-v�A�u���O��M���޻�x@���b=p�`��\�
3��7�-�B�D��8�X5��M���u2���P��z�NȰ�f;�3�2���p�=����&�;��C��
mŞ�Dy�Bެ�eAj����Lo�9��_8ô����ߨپ7��uf�]m����������β&�|2�v�"��"���ņ�ؤ���kXW��jݕ����@�dç�r���$B�[쐏�:A�t��=ҝ���B���D9"ipmH`��\�V;.���څa��(D�$�i����ò�NJF���Ĉ�pu�Gx*y�di��۲��CR#�m��㌉b�E��-���Қ6�U�u.N���,;0���\�snr3�W�ݏp��6�OG��@��	)xH��E���r�ֶX\ǬZkF_�
�B���]=R��xbd�8hH�i�/R�9|1�S���G�MZ�ߍK�UQ	q��"cӧbo��o�+2�g 	�3�e}P_ Pp�\�\� ���a��9O�
�����MB��T@znj������ë-zRؔ��u�8�֮�Wm�ۜ@��y��\�g���ˎ��$��:9����	c��Mk�t4�Ȝ�V�6�ц�M3n/��jt�m�A�}�^&S��1E݉�
6��R�2bV���\�
S�$�d���D�ڪ�k�!o�޿G��e�O���Q3��tR!	�V��&�����$?ͩ�ȿ�$�k�A���c��T}��{�k}o7��]1ۭ��Hӧ�e+*��e�s9��~��Y{�������P4�$L.�����>1����QQ��wG(���M[�o����
����������m�8�y�m���<�س��CS���N,�|~�M��.����
]�����&�ܡ5�,�5�2�^���Ѷ����Wϳ'�>x���U�l!�ܛG^���Ѓ��.
��*�#��E ����x�R�ˋ�C�T���N���]C�aͬ셲R/e�Q�_EVZ����k}��������о���(k�-�b�V�@y��ܤ�P�~'$��ڶ'���{���Sು��Q�E�۽ZA��Zq��Z���p!��k��b��� 	��L�1�p���iYb/~*渟H!#r�Fv�(���E� �/�f�m_���[s�c��A��  ~R�A�����n�ç��MY��(��^o�J�B�	���M[�~��^J�u���O:j�I�TפZ7��&ƥ��Ĺ��'��KK�ڏ���-C��-_M�D ��b�z����$�!�n���`�IKs�UjՄ�� ?G�-*�|�<X7�9�Ͳ�س^<���X�	�n�4�	�[�m�Bn5�x��0-��<�{���P�u�����^ϼU��Sﳆkީ3۫,���X|]-��x��h���z̝?-o�	r����5��U���K��hp�3y6���5��A(*�&�L�25�r�"Up$����ɭ�#�@@,�p"�rx�9��Wp+��e��1��55snq�+��3g�E�8:M�C"g��B���Ǯ6�ᵼ�o�*�b�-��tͥ0d�L/a���z$��6x�-qlc���ePm�
���֙eYU�Ehj@ۣ�ɲ��Ԇ��!�eLa�WA|��S�!��<jla�cX�qP��+2�]ӓ�5�����j}bϓDD��ONEf�[U%��?.1��Cj�X� ��ກ���]S���nG�5�z���[.7�]�˄��lj�5���j�Et�ڔ�3��?J��9A��i�6n���,���,���z�-B�({�5M��O���`�T��=fVƵ�9������%��$��Y8ª�O7�����Et{GR�3�V��.��Z�A�˭u�4���-���m[tTђ�;�^�x.��2d��#���� [������8@�C�1�)��m�`��$� Ѯ5����7�7 K�ĹXj���w&	���w���Z�8����!�|�'-p��(U�����;����SC=�I!T��$���y�cM����j�(|1��G���ܑa�H��SJR����35�����v�X��اZ5Y�e��m*2 ��Q��Ö�b;8��"�w���X�*-*P�o�t�!�*A.<̱F���̗?r�4�O�)�s�����y��aAʮ����Q+*f���!�I�I���9l�ĺ�����3t�^'��.p�_���W�%#g�0{!��������c0�,��!� E�9v�N�{f�řY�G�BH�'"E��&5�㒛Q��,��ti��f}Vf���J��53x�{Y�w�w�J�F"9
��~²,�n�\�s7�̛ie�D�o?�a�@�01�l��J@���=!^<�{��ˣ>zm��T�i�h��"T=�Fd�to�M�nG0ka{��^K2��F��>���CmoB��灷�:>�"��ր�sf��Q�Q��r���I���o�܃�zAA�O�   k3B�n��3�a���0�#JLQ�gI��F�Ė�X�oOb�D4:v�~x1��Ȼ�oQ	Pn-�P;�ѹ{���oN�g�L�}�L3��G�j���$�~�:hO��G�~|��F¬Ps|}�o����E��W �؛�#��P�D�V�9�-̋-Y�f*����r���ZDJ�Bq���}]�鵓��>1�̶�{*�zR4u��t�Eƌ΅��Hl�<	�������y��'�v$�||�၈���n_�4�:�gB�tUf8!!;��s(���/z%8�.#�hq�W2��}R�6��|��\+@��葤Л�%�����e�fw��)�6F_l�h^0��S�S�$��F�f4޵�|�^`7�[+0�$F>ߤY�[�)p^����㭀Y�-+���"LW�`yw��uMDU��am�x������ݦ�-�G�5�[j����$�F��:�B �x��hۮ��<�l��"r�V�E�	�i����No�Sܲ�94a�w�2�K�dfLa)9���5~�QJ<��㎌9���R?QZL(�C3�Һaf�]_�M�mR�C�ǚ�a,uC 6Rm̀s~V�m�6m��r��Q����0ޛ~*N�ͻ�g|Q�C���@»��y:�tS���֩�/[���&��F���{{�/��^���[��ԇ����x˧�Lkp&��h�c?�&���U�1��7[ի�����@nކ�[��>����.�~Ɣ�Z�^���M��L$�@���H��E�����A�:��(��&4j�0H8&��V�<k��߅&V�<7�%�OS�3�IL��q�Т{��گ|�h��;���FF�+�A�><�:�3LO��M{��+�/X oW�X=���GȺ`�xU&��?ƩrXǑ��ۜ����b͡����.A��ٗ���Q��x�Ug���:/�~p�x=�{���ͺM��"1�ό�$��O-Ը����r\�٭R�\M$͛Ϛ�/�������N�D,���9��3���s.��a.e$�b�KS�E��Ú�=�Jψ%��qr�/M_2'e&۾ɫ��f!�l�3�X�qW�,)�)�#�;S�b8�{fB�|�G�ٞ���$���惨Z.�o�v�-H\��ipU�:�Gf��:X���쏠h[�`_@Tx�f"��Zr`�V�/O�������{��s�ʒjQ����'!�-meN��T���Z+?u���%vі�mZ(�N�&��S�|߀Lʳ~��֢��מ������&�IYX����*�״:�?Ѓ�����l�SM��,�R��{"�Z�U?���1Π�!a�^�4>�^{�f�����p�&0�G�܉l
�<�����j
�� <hq���|ҞH��l�Rܢ8����%�IZw"į1����Ţ�¬2ܺ�P�V*�,৿�g~D,�^����u�ڿ��6�KL+���h z ]c�O(�]���P�G�4���z��U����P��Y�8�rD�'\�:��S��w�/u��[Vy4c��k�<��b�(�]��@��R�x�cV�������*��@t��$i^�*��EI�h!��yH_+�+i��ݍ#�Q/�J�E��H�N���_Ji�s\� �FU�V��R�ڒ��}�*��7��'���TԾ�8�a�g��ֲ���?��)a�ك-bi�2v|R3��gr�z���,����j�K�t���c]�}n��!��_V)�78�*�"S����:*����Y�����V�*G_!jtRJ�.�t���8��F��H�l̯$�H�ŻB�DTጭ6��:H���'�QLWϚig��P������I|O��FN��4dnc]X����
��
r�Z��d-]��6yvM�E�H�W&_�g�n�M��\sp	�Qٛ�@� �7�Q��G��Y�;K�em�PA��|�J��K8d�U�Zz��z`c��=��0d� �"	nif���lQ� Q1�(�Ț*����vԉ���}&9�l�1l�T��Wuy�wT雲��BzqC@ƾ�^�ś
D|p��!)�\f2+B�*|_��f�������٘��?[����I�w����y������ �q�4����9�*?C�Y:���"�;����bh�1B!2��S\������B˽YL|�HQ#�����b)0e����ۧ>ׂאu�ZZ��j.z�,�`Wt�֠���\�S����ۛ&�_�V A���ۧ�¢;��~|��`]�
�R1\��r @ը&u��0
)ElN�i�6��>�f�&�'2$##��>���h'P�$E ��+T�8�.��s���ޔJ���6 GK9ۯ<�zbB�}����8��R�0��gk6	IN��6&�]�H�:�X=��f�{���w7��.�l'����`�qi'n.�kV�M�����#�@K�� ]��K_�9R���P]Hϝr�^	��CL)q�~�
:'�z���t%/)^:n�jQ�Ҵ�{q�oTz��U�O�0�759C��r����X｡��(a�q��N���3�0�@:,����mav�Eܼ~���PN]"|ǡ�tD����?��@T�gha�;��l�9�"����ZѲ8X�	�r�.��Y�����u��!��7�|��S��@=�Ɠ�Z?��1���J��I_e0w���i{�-ia�ǵ�Qu�P�{��?��s)wI]�h> 9������^h&B��>�S�֦dxa@�@�K��o�����-V-�B��g�(�������X^!�����=���W@�� J; �r;"�8�q��^�K�cyu��/"0�i	�!��T�