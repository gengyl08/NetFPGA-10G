XlxV64EB    53dd    1130<l��6�w��e^�EXӢ6�L�<P;!-S{#�;uA�Ms�k:�X��_��4�W&#��.�l���dL��B�IϤbjj� �!��U�zҶ�nd=�xLj�?C0[>����~�8��j��EC���r5�I��ݱ�mD�蚿<��X(qY����D*�ϓ�Ng�$�ɘ��7�zږ�K; �ncٓP�7?����77֖�:rW�v���e<�6�EM�o�R4�xl�W�n�z[�/ ���xG�q/>hwN�T�뉍�fʹ�cpU��V�Yv	M�Q̺�L.{F#(~s�Z��q�� �([�<!m\r��J�����\��Myj����c��BQ�7W���I��&��
���E�JaV�fJ�#?%F`ޔ*��;K���G�4�N��M< 鉦M�u�3$�+�7���r9�����Y�9���b��A*�j��?hx\���	6TM��-�/���.�*����.a�G��xsMa�[{��`���O��;��u�D�d,�Ni� a�.��U�����g�/Dy���k�׼a���6�x���BW��p��e��	�J}��# 9��Ёmq���M򀟼��vո!lP>	aT��x@�8�N%���N����j+�������;������R<k�(��/�D���i�."� i��W�E� � n�&!DZ$z�rםLq$1m�!�[7��ǽ�D��[�ؽ���@��Om��킅��A�\�2����0b�M����n�fTw���GE�T��+�Fdc4'���rט�y�6�ʉ�w�S����)_T��	bU�c����`bD�����,o_t^��>gל���K���6·�O�����ߍ7dЌp�C?oA���t�	/ �l6���RA{�j]�4�@#'�e��m�8���V���E_�̤֌ը[(��Ɉ|�P:r8Y؎׋{|Z��^V�(ђG>$N��g�s�_
��K��	���/���aK���[�����E`I�����diY��d!�&K��˃T|*Z��ʤ���?�	����i��|�#�Mg������@P�����ҥ�ئ-��l��K>t���֛QY�t�s�ԗ�V�
EG�1���`�"�D�t��G
FZ�Q\[� c�[����h�& #b��j
���r��1-�����S�k}�܃�Hk@�1�� E��7h�\:��8�����I���y�{��FJ�fvps�O�K�%���_q_3��ũ�9�b��T��[����#ɹ��c�ְs�����+A�}���5�Ӈ�/L��Z����G�y��B�M맮�q�"&,��>~���b/V{�; Vj|���2�!cZrez��M ���
`���ۑf{kYq)-2?�7�"�CI�N�ڱ&B�A�ں���!%]�*��.D��|�}�H�t��vgҐJ�#��>��k�Ƞ�4�k4}K�#	�r���|�\��4;�7�ƮWZ��>C��43{���ma�˗@wqDh��.���YY�|�e�9�[A�tZ���T�'!ݯd��dw��+���4tO=�;�QZ��x�h��[ZH��|�(oͱ�w
��*�m�LC}ȍ|�>�g�d�_З�����=1�h����Rl�m�C��۩����������+����f�G�v3sqعo�.Ub����i�8�XK�욻��Q�R���ã-Ν?5��
��3��<-�����=sj}K%�[�Ȉ�����P����X�^.9|o�����az���%^�p3�U���kIy�6}�L�����Y�*Ef��ω�;0<�g�����K~�>H_��0�5�?4���'�o�6��- ��e+�.���(�>����|�2�+1����&��w1�w���%\7^��UK��dR�he�K�Z;����ѐs�ƒ�`��Ak,�c(��?�V��S+�>���J���2�F3..��A�ײ`
z�t�K�&�K]�K*�^IH���u��jj�̜����oI8d���S�U/�ݢ�b����o?2Iy��`Ilez!_{Te|*�h֦!?�Lxm����F	�:��V�n�1yX�юЯU�\��&����Ďo���G�x����UA� ���8�̷���CV]d�%�L���e�6]�(k6vN=��TB�B��B2�s7�`�w���C$ �`��9�QWm�z������>^�r�ϟ.���g!R�w����{ V�v'�F������#8�����HͲ���5&�!��V�fw�J
{����,�[o��aCA>�q�� ��u��)%��g����M�?��A��5߳����C�4D�q<�h�BM�B��u��y�U��j���dSp��8L����Ryh�Z-U��24e)Y+����;F��î�{�S�K�V��rt'Q���mf.Xg���5Z0�ȇ��ۯ����0R>IHID�&,�r��O��� f/k�"�c�}����J�¢�a:_�RW[����Y�WoAj���ꇍ��+@69������t����ή�y�%�1o�v�{@ߵr�bߦ�_�,���#��"t�$~ȫ��6D�\-l�Ե���ڃMp,�'��c��0�C�An_T��V����C0R�����X��xM5�P��U���@�ux��sn�?�AS�����_��(ޣ\e���)q����(GzV�!G!�_�g�.?M��_"�vK�*��U�/|��I�u@���_�6�����r��b@�ZDf�6E��uA��35j�<|�o��/�p�Y� �G�&�%>9C����T��f��e��B�v �D�٧����<挚�9@s�U���9wô���>k��r"�O
u�6�]h,w@r�t�+W�)໅yO�g��C�;a��>lFs��\j>B�BԂ����Uڄ'k�r@F!β�d*��	0�9@�h5"�2%��3�=����#�23Gn�~OF��>�D�[���=�|RZbА���%"�Ǉ��G�h]o5DA�/a7�ʷgJp�8U�b�#�M�����O�]�gs<���x��o���j�j���(*����7��o
ԴRD2&`b��)��POo�{��Hx�7SGqC�Ώ����UA�Vj\l�ߞ����z��P}1�|%"�wP#@S�Z�< U�������V�x]�N�6A2_.�;��El7�a@��Lu��~�}ö�o����+H���.��Eu��1��w:�}Y��[~�L���g��.��n�i*�VR���$�$���X�W�:3��JU�n3�E�t\@ݜ\㱄�h�$�����T^\���Jpv6b�:C�]?�K_dz�2EW��7M���L0q6x�ls����e0����}nϡ~s"}x>�^�Q�����_�ﵝ*��`ψeX��z�/�	�_��Y:�BZ�`�7��x���GD�xO=��|��*�l��I��u�ȃZ����Z��Y��Q�~�`���8,�D��%P�����T?'�!���[t�4�T������)��]��9ӳ�*$�U�&��A�­�02b�%!�6]a�B�4���ӻ@jφ1�������>p*yI�b�"T{
�IG��֙QV�#w�-�/��XR�/*R���$)v�@��p#�Mmտpd����=����h�
��^�$�ˬ�?x�*�}��������mΎ�L-2��V���ܕ�L�k����]K#��Txb&�m`a"UD�shh=F)���{��k�W�{�S%U���)���-vnp��b�����V��D�yF+R�O5���Ɗ��rͳ�4p��1$T�L�&�"�)��8.��������z<ux@c-4��'��)~�j���_Ӏ�y�uq��_
h>t��X���~݋���s�TSNױ�ݓ�Dzs_F�1��Y�2�z�e��q1U�y�F��[zR
bϼ�UX�v�.��ؤ�	�ϼ�JN����3������19��J���8���(�Y���	��N@Px�QMbc�`�]U~S�ɟӝ�x�0���C%/t\K�P��ҹt��߰ii�1�l��Xe����BMRc�7��d0��ۑ��D@�	�HY�g�(�%���?m�OH�|���ml'C�~�S!Ox��#�(u�H�+���`#"�j���˷_ПS�h{%�D�W�p�}��h$���&�����хݎo�M������������!���H�;��� yC,!˗N�zw��
d��l������쩓��2 !wu�� ѳ?Z{B �Ѻ�ڟJ�8SX��A|�¦e)R6�v��X9N�:�+AG��EZV���\�no5��;o�3��N����DYux*�#-~E�