XlxV64EB    584c    1340g�L1ZɓrG�%�t^���64�������v��3�.~4��U05U۸kg��`&�,嶎����[�}�-�b�6�%�u�M�	�d]�����gb����`{,�gk��^n�!�0Dtq��/�T�a^��_��|��{?�f��R�1�����f!7ݎ�����̿ �/��ژ�C�meX�ޢ��->+����`4�����C��G)�1�^��wb��K'-qk�-��(xmc7(7��o�ޚ���� �?H>i��Aš�%�>U�Qa�*!(I��gjn4�+P���p�M8߉@9�zqf�E�OIj�:ѣ��`TGmѯ�4�`���曣̍B�NH�1��P�k喱��&�")��s8�F-mHT��#�w
�͛n��O�xn�!��QÂ�#�*���C�|4t=)Qb2��|;8&&c��S����x���W��z���BA���Y#�E��?����.Y`.� �w��	�~�_!e����+gF��Lc �����iB�c��<y��Rb�o6���T{�;긒���]���{?�ߙ+��qtT�-��6�_�ˉ�j�+���͗����]�j$��}�V���_g�M�@L��e�&������^9�)]+�gތ׽;6֍�_���yEK*?�um�
�~V�[u3;&��M��S�S%>���Xd�l�a9���(��h�yՊ����Nz~����9�	�P$�S6z$x19��KW��K�O]J�.IX��9K��؈�l~{
���P(��`�}&���v�Fr#�2m��
ȩW�Vܿ��kc+�UBl(�cI����#2�݈p�b?�-����H-x�w����s�Z��u����{������D�J8��wPi��(.�
M~׫W��@�q�JE`��y������`��X�o�j�r��;
?�z\<h7���gg�[��g��N�*K�r���U��3����r>�q��=:�V䀻i��Jr�Y/2�ԅ9V���s�)ڸ7s��,.H���/�;y��Vz���|�O� ����񖁽���*p��v�\�b��g.�M�D�k9�h-���R����i�>�)-Z	^�A��%��7�����0TG��g=�n���d�I�/?�P���tA6�����h���г�~�ʾB�7�B��l����5�@�m�y#8�Jy�Ym�ٜgF$��/����U�����N����ǥ�-�bm��A7+�s��|��Ư�Ppۖ_�ZU^e��9�#�Ak����Q���W!��+��1&o�?��.B��n���c���X���>���=ķq�!#kobʉ��E� �<�)�f"��chGLA�W
n#��-ؙE���Mߵy#��"I��f
�0�l���\#i+��ۃX�:��#r�ׂ"���Wͷm���~x@T����N� !u�45r(Ϡf��� ���
FT[Z�l�|HLGX�k^�r��"�3u|H��'���e>�s�:�L�N0�]�#O�<��LiB>ڊ�SVo��R��ZLK&}�V�"�n��'�M�w�h��e���5}���S�~»R��7e��������53��]!)A�����#���dc~��h�B.�@�pF��B7����B|�y_P���W�<�cc*�H6�#\Vk��<��NE���ϦI'���҂r;�t�=ٗ�u��2����E&�%����PRZ�'ոmy��W Q��X�Q( Ш:j{�&�L1���vlP!�c�D)��I���w�4
.�ZFǢ˫��$*��L�	*Lw�Ҋ!��s��C�tց�0c���}d���X��/��/�y5���ԑ9����	p�� �'y���P�U!��/�z�S�)Ectp�D����|5�Ɵ��wI�h�V�����"4��ђ!���_'�>��'h�@��Q)�O�ƶ]����"�7r��IgHC�����d�wtAP��D���î�C2A�n��d��6C��$� ��Y~0ѽ| �)���M�WR�e�yǼ#､��?���Ė��c��
��?P�%Z!���33��b��dP�Y�M�F�48�7��'����V�:~�����3.�a�:H˥��X�c�PCX��`���q�&���?S�g�?���"�w��I:��u2Xg�^tm��mh�|HP�t���L8������j�u�R-��zX�Ϡ��g��qV���v̥��k��!j�������־D����T����1"എ�ga��!;h����n���� #��}����Ws^���e��״o],
���r�wό�EH�^�\�)Z7���LF�|m.�ە�I*(Uu?�z6W��Xko��!o�U��O�WƐ����e��Zeb��ؠ)�f����z���ȼ1iJ�]S�^����/��f��oo+�}�a�"`u��L.Z?>.k��8C)/��4��ώ^-��^�Ɉ�C���y�A&�s}����q(J�s/�<�c$^W�7v�σkue1w
�MڻnoE��@Kf 4Φ)<�Mp���*���(�j�C�=N��/��~I�A��l
A�����g���{h��D�K��9�6?�y�n4���#�:?��ج��E-�83�F���: �K��s�ãG�8�0���X��2�U�U8^F��А<J�)���P�<׋��� ���.��Wj�Nu$<Q�pm̒1��^�?�+6c��Y^3v1MC2w��Ho!BVb�D��t���xzV��Y�p�͒`���V�B=�r=����Cp����[�&��v����9���8g^QDy���+�[�L&\!�'Uaҝea3�ĉ�Ѧ|:�w�#P`��$ۖL�d�[r�te]#��sj�9�N�2a`�@{?���,���h�{����Gx�Q�\�9wp�o��3�r��C�h���P����U�aӟ9l��ۇ�Qm�[����B��FG���ݞ���W=��Yb�zk�(�s�@�wDЀ���o�����hc���Br�HW��i����aħ��&F�y��Z����
. �56}e"�;
%�Y�P���6\�/����t��CuEެ��u�m��!I����ݹ�VT}��h�8�{�2�G�+�4�2���+�{7JR`��P�O��n�4��������㾒�����tZ��� љ����?T�<��tQpET�H��l���*޼�\�`A|x��j��m�oHe�,�3���.X��Z�
�.�j��@�qM��Lŷ�-����n���W4)��mF�	�a�(l��H�'�ڌ�I�m�Md�ŵw~����UM�u��a�	���o��q��D���תԛ�a$6�R`'�|���N悼������j�
ႆ�^�U�\,�Gg0��ƿ<���rp�#�ĭ��Y �)������A���2��T��ӃzO7�m�P5��]���0���<�]�G�W�f�Q��ϥ]���H�΢Lϖ�,��5}�r �������K�bv�K-����7��MJg�.��y���)w[��Z+G)�!b��Kf"�׫K��+�p�����5n�@�S��2=Y�Κ���2�l([�6���x����fSl5)�>w��+�B�޻V��$M� Vi��fت�g�u��a<b�@f��0Uû	�����Ҕ8ټ5G����|��"��=f��&����\m���r-oé��XB��qKG��#Y�EY>���p������\]�`����N	�ܢ̭�m��h{��3���}!EU���I�z<�#>Qܳ��&�__��b��c8ѓ��l���gY���$A;�y�H�ʹ.��Zl���d.�Մ�<?WMy�U���F�%�r!XS�F�5��,"��>�~����E%/Q�`b�W����8E��3����U	�l��o[�����!ʉ�HՄ*�wjCI�s �K���wF��k��������%i��O�]�у�I� ��y�z=�r[7�5���p��J�c��RS��Q��/r�^"�}�J8I7,�Q7�9Mφ��B�A_�]M�$PE��� T��&��UTY�5���ME�؛̺$稥����-��WN�47����8G���	����l��j��L����(�`����4B{I�	\�_�!2
_��Rf�rÕ_�l�f�����m����&m0#�5�4_�B
�-�_\4z'���19���by������y����7If><��~�w�%%��O�j��O�f�dq����������<	\�kU\�n�QT�hE0|38�=�hJ�c�$�.g�E���+���� ��M����|᷍�:�hKN�G�z#�1
�Ѡh*d���eEƱ�%�� 5̺W�	��G!�_�\�B����ׯ%՗�,F��<r+vOyK^��l�Y�|���Xm��3�����rh<�u���֏p���G�6%+N����g�������-�<^J��G�����S��;4�������9w���xx�*����UDz����]h���KA3���YG�����
�����[�Q&:��}X��6�wu��N�
�~�R{��#����m��],�m	7�rW�*����j��-I���B$^���LUO�oe�D����d�m���e�S� ��a��~1h��S�gb�m)}��L��������UvnM�ד��tQ/�˼� �e�&Cx�VIq6\,���n���zz.$�t4�`��O'�d�P�R,��bX��&��$ʪB%���z^-okm-�f���t?��UrD��j �u���TZ@��r?ٔ�F5�E�mB*�Z	R�,��Lpu;��e��JC���$���xTD�q�;�]��P�A�j��~�s=�;mm������qн@P���^�6~��N"G���>p�:�
�^P���W�� � (�%�t��pz��dEL���