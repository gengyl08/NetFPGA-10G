XlxV64EB    31f9     dd0X	/���Hl0h=d<zw�#� ��N�g�0JpO�gh��֭�q�+nQg|���%�2��!O���0�I����#��6��ck���_|��"o��?I��74�/)�˺����Y����<�+�7�RZO=$n�h����:��Mƺ�-&v;�:qrL�?�_�
cbHH|C�� �
Bߠ&��%�0}Z�DmES��ν���Qf�e��iǻ
�	����9��LR)�ע�B)�⮘%���[��!�����nT��'���%M8cs9���Ic���Y3#��o���I$^�i^Sm�.؆57��߸q*
H�a�F�$4��I9�8r5z���Xg���W�+ؒb��P8�es֐[���>] t��rm�����ۯK��z�$�[�?�mV���ٔ��6	��e�2��w�Մ�v��A�|^���k9�W�kƈTS�s<�H�T��v���,c������>�&]ʒDT7����#��X՗tH"
�u|��W��[�A��M4�� ���|1R#��\�z���򻮰<P$� �sG�B%P����$�5�����+V���R(�W���Z�<D��on�� 5�kA�t� �W����!��j��$����h�&�}��z7��ͅ�޵�����q�g,F�/-����y:���`�}N��� �
s#R�T
2"B�n�&ڇ��V�ĎV+M���z���kxM�	���{!T�˸.'�ߺ�٪8v?�"W�����$$:f���g�O�u���]���h��+���j����@�!w�yv�S�v�#��sC����Q4������̹������M���<��B�S�;��sc��H����$����Ah�A
�.  e�G�gA�6� ./�3f���QIu�Q�!R��v�G�2>6��8��g߄vз��>���m�(�ǖx���k(�T� �j�5Oi(��߽X�p�)k��V�S�ؔV�vU�n�ާrx�����^�(ؕ���v�<㠳۾@�%�>�x ���S�ʟ���؎��|��^�
c��C�63�����
:L�Ko�g!��F%���5��n���i�4���(�_Ђ���4��j���6�Ii�h�O�G:�䕪U�)��w>�G����AuG�,x���A백�F3΅���ASYR\���N��c��:�KBc)�R,����;Wm�:�O��L����H� ��!�.z���As����oq���!�� l(z��Y��ܦW���$�`Љ�/P���B�����9��F�:������%�s>�XV����v
xC��l��9z�dj�0�����sT��
ߒҒ��4��uL�ZQ�o����x�!u�Զ%�����#tK��r�#�S��J�^�3P����Z��J����}��kV��{��&r���V�b���]be�A0O��^����O��+���l������{�AF���C���쥞zi5�M�/_t��K��0~]��w�g�(�=�׹�~���(g� ��g|۰��t�5�py�%@�j����`w�qw����~ֈI2��GC��\��o
�f�#:��������ob'M���DE0�9�\���'l>׶Q�"Q48����k^L���-����[��f�a��d�DH��2��ЋMb��x�up�R�}���Ќ���tD�o�x^ޡ>A�?�d%�8c\�8�E��'���Ci�G��f��☝s��t<����w�٪�n?�5��a����`kfj��;$���_9�W��݃����lUu� �f"��N��u��1R��?s.6�u��'婍C����:u��}���Z��"�_*$���sT������Sm`�r>���Б��ɼ�����\2V)�y�<<N;�=�e�˾>��di���JM7[��캿�K�;"�ؠ9C-�C6I8����Ԓ�WO~^���Y] �4m:h��e�Kѽ;E��8�!m~�r��)ǟ�3�_h��&��4���;�� z��Е��NDS�:�(l�Y�Z��Z��p�B����;䯸_V��bb��s�?��|��j1� ��w^T��/���x�Z>��E���A)�'�1��
6�����{x}�p�^%/�k[������W5K�3�~�:�@z|:�
x�
��;��v.?�:<��W���+�^4L��pl����t����
K�G�Y�]����}���|��j7s�<���'��XG�`���%ƍ�3]k��G��C ��dUW��(�%@�RF�Gy�ވ쑀t����vlD.{M߳�����}G5Β �&o��XG����EH��o��x�=�1�k�ƤhtF���L��'�^��8�S���صFBS�3�x��](k� �KSB�T|A��:�^"��@�2'3x�߅
�,̓W���S���}F��۠�j!Z�4��pD�.��|hU{���h\���yx�(e6Xj�{�½�	s�.`�O�^h�Q�>�[��HG��L:|���� ߍ�|KYtK������'�<&L���εtþ/����V�����Fx��g��O��6e�ѽ��ע|�{SY�}P�x�r�s�<�G�Q�bIX-*�,*�\'{

�J�92�
��'��̭�4gZ���ݴ#���F�<����M�����]�I�:|���v�_�V�ѷ(�R�Gˮ)�D��!>���.7O*f-^Tp{yy�ң��!h��&�Js�ࡒ��`�~��踒iIY��k)�o��:-�9�>&KA���|;�#�4r�-K�W�����]����j;�6�E»7�jN�^8��^	�u3�έ�$qⰏ4���k�2�:@�0T3t*�{�5��i$�aX�ɵ�e�����_��F����l�Kj�`�7aE@j�T�*z)qY��%�ku��Nki/�q���g�����;ҧ��NصIT�n���K��/�ժ[)U��M��>eb��O�x�ޟ�U��/�t�j@ԛTybx�^&� ��n��g�'n=Sz�-����k%W0��a�)�M�r1J�5�;��C0��Ǆ4aK��v�2vD��9�9j��<z�p]I9��^,���'�����J=���6��������b۔�<�i�Ԧ�<��੟oF�Y~?���"Ë�#��A��x���+f_���G���T�j|B�f�lJ`�w��=���Os�ӗ�D8#X�t�S�?�ͭ�A�r
dhpp�6Ԑ���߭7�~ɕ��suAzu���c�?��������
f.�Hդ����}�/���:r�*L��JX`
\���c���t���f*�4>���|؎)�q���M{U:;����7p>�S�m������m�ė������f�$#9�= ��A�lU<~����Ǆ��5n�u¥>7{t%�ŉ�=����[ W��Q��o9q���:��I_'c���D�бb��0�:�?eGpR�Ia������R&��]B��"ZD�I��