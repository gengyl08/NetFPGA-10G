XlxV64EB    55d2    12e0���A�),l��P�M��a
+D:I�����=S���%�N[�Q�������n�B�Ϙ�#�����.�O���\2��}�#�YJ��*?Ŵ����Ԡw��
�hCk�D��j�7���y��H���7��ѥ+Ͳ�� �5���޳w�x��Z�Y����
�PA�"8i?<���O�@�����X(X���lK�K4�)���UܪZ�i�^�E�����cg2��
�?���-x�Y��Y`m��� a�z�O޳.PV(�s<���#^���/�?"���A��xH$�:�qm�{C!.�=a��mhMt�ء����&��l�)�J�V'H���E̾�ġ�(���.�X��	�R"��<�"*L�p6gA����q�!�u7ehn��爛y������c4[�1e� i/Fv�]JR����e��p���	�n����ZH�6׈Z�_�x��ǝ�%L��y���p��L�;�7�0\��6���MC��M����(��\��v��y2��ʀio �J���ZQ/��0dҕ�R�����xڟ�^ED�A�7�4������u��l>��m��D�}���ӯ9�N:�_4�_Ye
 ��eq�!�FH�[8g��Ѡ���i~�(.��֧���j���~��;�� �_ZWTp�����/��8k��1]�D����R-̟�f�����Z��l�o���S $��D<����,�}�?�*
����U��wsl�l4ن�R^
��IӘU��5$hWF$N�'}�~���'�v�N�٥#Ts�"�����p��Ձ׾y�p{(�	�N���^��ŏ��V�4�EŚ�K�AY�/�����������䣪'�N�~���&�2T�[��M� �x/	�`�v� 21���cGd��<�Ćj�p�s]�N�x�`�:�7��.��m�ej���dg[�M���6��?>��"�@�#����E�+U|�X�a�P��+ɭ�B��[fXu��Qk�
�V]��t�<�����nJ�bw�j��f��5�e Rr�u���g�raT��⯀����3�~���E?۸�W���Y�夔ZD�`18�KlR�Wy����>XC���b/Y��n�\Ĝ.2v�+�D �n��ޛ㍱
��EZ�Ov:O,�)E�����w�ng���
h�{�z�Xm@��R��l��B��ߙ|�[[렎q�O�)��>`��a<@�H� x��c`_��l��
��t�ltҸW�oE��8ϛ�E`��st ut�1�D�#��g�#)�� �jߝ���4.\� Մ�[�"������l$�b��x �����~�q�z)=��q�[�JY�0�<��*
Xٝ(g�6Tj���&�\�<6c��g�Mq�r�����L��K�_o�`]hȁk�����P^FI89�I����ʂ� %<yr�$�����J�_d�r\ߣΚ���_�˔"J��f�7����Y�����vl�x�~Ô�C؋	����I9Wֱ�޻���)v#W*��h��j�h�o*q%�J����򪳳v���;��6��:dK��fӖTLb�#0�%�caq-��Px�Y���>�����V��0=c5*n���~�Z�`b7��+W�q7�o�a8��y��	6U̇Hc�՗��s��ܽ��/�V���/F���K����g��)x�R�w4ӄH���>~sL��/�0,l�S��s���E����#>�}���Uu� �*0%},���E1�*́C
�D+!�Im��Q!��s�$�r��d����qXy�FB��\���G�Z��{�s�B���$�/&le��Y-�N�\���XK��k�\չH@�����J+V ��nV�Hu>�O�T����4|�Q'"�g �M;�~�g���k����m�lUU>�s��kb���.�����p�}�h�3U�G�ɓ̮@*:Z��q	� ;MyT�6��}$�3�c�',ҽ'Ψ�����c���k�:U��"LV�Z�א_ 't?�Ǒ���<��D3��*�c�Vj��i�ѭ��.dY��<*��A90%�� 9�$�3�Eq:�
ПäV��Ь�Y�xȾ��8��E�����h�MOb(|D�H��"V���]ە㉝�iͯ���p�T�M�q��L�b͙'��{\���xDmb|�;Gj�#T\z�l��8�;]`OO�0�����@�r,��
�CKT_'�5RKR��T}"P���z4�H��8�'��8<1Uw�����b�<�Z���R�Z������#kL
�����<5�~�	�l���C\7��0<���]�L������?	�-����.��gy��`�����<���\�}���iLm��sA9�k��s� �vF"6��A�װ���x�`����xB�Om6�6B��R'�i�������M ��)=Y���;~��"q�������<�V��dT���NF�����B	t�s������ק��$cA��W~	��g�(`�QŞ�0?{��*1�D�r��2��^ܠ�Yv���~bU�{�C�L�ƹ�K�P�/A[`Nk�i �\�X~>�������+�;�f����c�ut� �K���d���t&xE�a�2ެ���i�T�<T��r��(�2)r}������q��c�RW."�)׬�մ\X4�G��M�E�q�@G�7���Q���*C����j�ybBT�Jˤ�4k�l���)#�R�1ܾ���)��*7nH���)� �M@�\g����lA-��IT�8p�&��a�c�xK�c1�C?ܱ��
V�Xg���|G޺��(L1��^�_X��Z���(Y��̙�B6)�h	����F���3l������>���M�!L��|>�w��Ӭ�&��;�(]������
�le��1���}/u�X-2^���e�)�n�d�9����Y��*:�~jѽتl�O'���	q��ؤS�\qg����🃧�ߋ�§ʣ3nH/7�c:�x�'lN�7Mi@ ��uu��?EL�f_<Q^"E��мy�'y��:{�Y`zw$s�p'y��Ͼ��{8�V�0�Zؾ�����0!���=j�L���w�����.���mn>���B��@���\u�WW)��>(�uy}ކ��e��#��/�Xm�ͺ�[�m�%��ڭp%��S�b�Q���r�A�^M��	��>B������ŕ,9��AzOX���Q�?Rv����e��;���'5��k���D{(x�{�U�D)
B���G!����5�͇uWƳHW�k#�)R<��W"�:
u�\��tD2~|�=��=��SP�Q��������|�T5�Rb7q@�II��2��n`�cA��̩�G|I!0X(��{C����6�z50/`}��ݩ��"�g��%fmS�C^����rumc��jk���"X�I⎛rR��wtx9�bA"Y�����~O��|�%�~Ij���X4�h#p��u�K<��$H9�N�y��O�}֭��=��v�a%��\(�T�on���y���$%U�mM1�q�-�h�ϰ�!7��8�o�n�e.��xy ?�\Nu�X��zsB/"�B)%�W�p���\n���{�JP|�^������~���G%�j�t��a(�#��k�}�$��Ǧ˻��T�z��
�i���t͵��`�Ȟ6�z�l�y'
\9��I��/�ƣ�Q�H�S�
�9����a�s�P������a��	zP�;`TE���Z	���R`��y��o��=h{2E*2iV1�0 �%�U�f��FoI�����Q�aA�ƕK5��|����$L<0u�����Eyԇrܻ���àۜ\V!����>������&�?���#�*�9h�i;2���D�45�T<��1��4y	�w��<������ޭ���4>�V��5��-ܼ���6:��a�U!p�fˤ�C���ؐ'D�9Z
5�I��i������"��k]���z���-���Lt��e(���!&j :;C���3X�aaUv����,+�<�ý��.�.���� �ގ��,����N��%}3y3�����~^�;4��1d�������R��R$�X����Z���ҕ�)�|�:�V�cz�;?��`�ƾ%��3M,���������ۓ����6���(ko��ԋ>��~T�� �ĝ���\�JK���t̥F���4:�)���Pzɜ�!�7>�mu��X�*�x�hQ&B4���ؼ|���Tx_�H�f�YnA��{w�����?6���\n��e��������m�֦�hG��y�m��ܬ�K�A�,��~&:��
�{*�ue��u�]��(2�E565kRp��N��'#e�1�+��a���\!*d/�Vطy%�:E��U�̟��^��V%n o�y�C�,`�K�~n���$�/X.��BT w������iQ�	�f`�zj�`�H9��e�W��K�^��)�0R�Vm�s�o<<9�����=�W=
��J�������pc�o`S�nV�h�$l�I��^W��c��q�j���~�8�"������x���#(�j:��&x�Z�w���z�U__�#<��A�y���_�!�:�%Zn$�y��o�$_j���<��%�H�vaZJ�Ӣ��N{�2���kd(jt����OO����w�;�V�ƕ3$Mɛs�ԉ/u+M�d�R4'8�51�6�(��H��d�faa��%:�~++�_�hB8�}{���HQe�>:�8���y��0�0�=���7�+س�A�)��P�