XlxV64EB    fa00    2ef0UpJ�h'��ȳ�0���q���c���y9�0%o�"X���pΓ��X <�T��E=��M	�߶�������蒋�I��c <_㨽~�}�Zʯ%�lU�&����B:�<�fo���pn�ڈ8�pϤd.��f�dv�bW�%|d7��Q��8P/^�3#���Ξ~R����x�!�%���F���6�C�)�j!�aP��b��J��5��(6�Q#!�l���O�Z�8���J���5gx�g��a�5l@�ݱq$��Y]e��2V"�=�+*=�
/���;��g1�� >=����U��둽W���X;9�3�_h�S�p��7qG��6ʺvqϑ��8��:iDH�f#�_�FBr��ܓ�!��C[����[���&V��u�Q����6���ŕ�[�� ��)���E���F#櫒A�e�FY�������U�b&CJ�v��ZuA�&��`����D���b���c�L�l�Ag����_�Ч}���U|�?�T/�r"��U��Щ�={݉��w[�Z�.6����g�� �������D���$�!;ˤ��Aҭk�1�d� ����LZ ��p]9�N������K��q��U�˭���B�u�͢Cri��U{�Z��cI`o�ۿ�v9Z�5�ȳ�h�LL@��=�C>Z��"��v"A�%�ߣK!rŌ@�0��\�nd{���C���۪f!�̄�vR��*U=��} d)d�G�W��t���^�S�U��L���c�������6<��/�b�3l����SX
դ)�F}li+D�b�$�GrSʻ�N�s��牫�I�8�c#��~bF!W��Aq�{����KĴ�U�D�W%�m�t8��$��^�д����g&������S6wzJG�)����>NS�ЇI'���-��Hכ:���|au-�u/ږwUۼ�͵�}���+�{g���(6�5#��t7] ��H����
R����gH]�d�~	:����R��`�{v]<��hi�3��"�cw�W��eqdHV�7<�����עj�^��IP�,f�����̓��N���q~mD��6.�����)�6B>5H�e�/`����\���묰�z�m�	���gU��N+fʎ`�g*�`���^���p�v�
�.Q�P���pꣲ�;���E��x�L����U�J?�߰�������!b[��S��r�e2��M��T?
>j��^�!df7.-���=�'-�9\�&W^�ms����֮���]t̠�ʦ�Y9`��ɒ��lo���Ҷ��2�O��D�X�݄?��%K��\|����w�6�f����"n���/�Wu�T���&�R���!�	�q�!(g{��/��j"�#g��o����o��d:�|�r^�|�����_h�r#',�]����H���NM�pt�X�0�Ճ�L�,cSҧ
� 0�E������Ϸ�g.�"l�;�[\�]�2���k��)-��[f�`�rnJ1�\�"�1�P�n�>�����>,l\��X׾[�#��|�����3�nM��T�
6��)�EX\�2�Ո�od����G�+��S4!��@$u<�F�+�GYR=&o�$*5Dk<G�k�(p�5,�ϮL�����)3���p~��pɫ�N���@?ٴF`�Z����wѩG�<f�I98����n��IE��_�%��<�x�v�� Ǝ9Pg/Iw�@�'��4)�_G�W��t F�Q��8y�P�g����	�N:�� ��pr����j�Ut�ga�8�Qvw#�-}�S��%q4#��`��[�\2����^�q�}�m��e�̋4�����5��<§T(���f�$8i����j!�،5�p��K��ڤ�@�c�W߅Ӂ���n��f1������6�v���}�t|ם��E;�%dmǣ�\�Q	)���;:rߝ����4Y��JT���-4��JU≕��c����z������ҽ�L��K��)^�d�`�:{�U��Y
�f(����)�m�R�\�6�u<�����7�m�R񩗴'��0���^�X�����`A|2H�[��!C�������>�^#�ksԢ���?DY��0��h�R:�5�x������"�c�a��,����C��������_�H�B�hRϓ�P�H5s]���k�+�,D�E��GCE<^H~�n��)�*����"@E��V|����:�i���;9��#<�Q�P㟟wr^�����>d7]�<�bC�#�r�j�pL�:�C4�okt�P�-*K�jfm�$�*��8����.]����4�A/���a�n>\CS���*u�Q�����9,u-�����v�%A.fɵN�+����J�%�,�T����_��%���?�ؑ1d�Wo�pU;M8�V��Cʿ�c�Iu7 s�9Ơ���(t�Z��W���[�-d���7��q�7!WY���/4�w4I1W����� I���fĖ݋;�G�Phҟ�}ȕ�؞5i�!���{B2�� �܃��s��ᶵģ/G��� �<�'Pψ������Û<z�Z	}#���y-�<�x	!a1�ӗh��>�+-�-�2��{<�DX��a�\��oy���j�z��AP�#�����(G�ܠ2 qt@9�wI3�q��z�ڬ�rX����]8�8�Ѩ�'j���+E�!��lN֡�(AL=�i8/|��i�����RKL�l�ԍ\6 ��>�R�D��R�ï�ㆉ`"Ӂ���ѓ5��v�h$�6
�:9p�w�
e>�\� ��ߦ�T�s�θ��[���<�(]>#F���x�~]����,@�?m��[i 6?�fq�h���t���I��k�9����2��o��y�Z�.��FYE�R�v�,��][�Ɠsi&�.����5֦Z����,�ċS�T�:�I���Cy+�@��4S�L;�b�C�!A��$�ɥ(����B[R�,օ�d��@]�,#5 0~�D�P�P��TB�`��=�=k���M��e�^sJgg1����ihX��{y`K���EG`1dj��' �!�s��f�3���Mo��e�H���q�Lw�}�j{�p>Y���kzH`�@O�RZ4Y�Tnr _s�@C�C��jΪ�����:M_�BExF#�̴���U��_��.�~6,3�Di�^�Q�i���:���A`D�h`P�ܙ�&��x5���"9এ�mf
f�մc��dr���K^s����ﴢ3	��M��&?3��ys6�:���ω������h`���S6J�+�e���K��L���<��3���KF{����&�
�� �QiO��+�
��m6��<�'�D��9E��8�3)���g�+\G��3#��Rpd��՘�J�l�F΀2u�dE���kY�=MD2!��6��q� Z�D�{n�9����c��Z"w��1e����m>��u g�]� .��Ze��7_�S�v��g,밟"�����f���s�x��j,��|�R�$qs\w���� �A5G���^d
V��kĭ�es��(ȍ��f23h �/\�.{���B"k��
[wX���(ox����K5�PQI%;��F��f�+��!���*��H����	�^�Z��A�ci�@�Z	�~7�:~�cW3���d�[�K���6�H�G�Roق�{<RA6&�J��!��G}�ܓ�L���3����	�FYIr�a�-�\_����r���ApS���<5�p�g�9r��4~��]fmV~�� ��n�d�7���&И�"����|2���m<�)���S���]� a��&��U[d=�X?}N���#�Ҹ�%�h
}����mx*�Ha�Ω��<X ���+ �#a��oW���2:,���h٨W9���b~���Wj�b������V��̢�W�C��۵Fk+"*�WT����htV��i�_��f ��Y7S��)V���nZ��u�I��Q�Ϲu��Ͱ��
72�	S��`�5,h	�<����$w���\
~-�{�Dj	(TD�����^�����"'�Z	�o��>X�N�N���Sg5fx��K�r�UF>�0tW�_�J�{��1W���z�YR�_166�;~���!ׂ�A	^&��/t8�?�����%�ҝ�6HV���uw2�G=^Km8�wn�C�H'	LA	.6��wZ�_h=���"�Ǒͭ,�q4ӷ��YؽUj�-�H�gM�ւ��'W5�5˯�@�������Q>�#�B�[HO%��E��ZpA�RÚ��8�jԩ�I�F���C�:x��	��<�Dta��/\E���2siP�w��{?�z��������sy�p~ ,�v)���AXW˻�i��1�7.៱��^!��,�u�
����^`P��Z,h���L)7�ǥ��:��&K���&k4���ʫ�]�n�����j�������������;LLӼ��1)+�5�)ߝ�����F���mw�4Mo͂B���h�3�}��uI�w'˶�zO�^l�;�g�gn'������J�B*�g5w�ߋ}S�xpU�ȧ�ĕ��6]όe���U`ft�_�����7�,H�n�!����>_9ve�A�BhĔrNO�%�`7z���dǻ{܋I�C��Qݨ���ᥳ��}^s�X?<K#�[A{�d5x*�xCs��,*�5ۭ ˼�e>����Ж5"8,�q�"M!Ū}��v���sW��*<�;�r��^�Æf<��0��mQ�>�g7��ʠ�Iⶇ���,�������7��j�,s��?2��i�<�m,cn����|�\��uO��� �c�/5�k�|��<}GJ"���a���Y��f��C�m�1f�Ly| o<7 F2�c�@<���TV���KrV=O�&QU78�XG����ݍڹ��꧀�e}`�!g2��P��N�7ō�����]�L�&��K�Y���z2�eނic{M���%׋��!�jO�Ѐ�T�;�����X�S��@������B���K)l����>«�T�C�R<����}�e`�Ry�}7�h��g[�Z��0<X24밼D`JM,�T���8H����+i���0�R�+��J�6*ʶM�����~�Zh3���p��bA}�r�L�2^j�6��� �P��� �-��'Se���Ô^2�{���zʀ��eߣm\(w�.W��&�1�6��t�|��{�[�Cv��6�6��n5}S�NÎ�2+�������_)ʡ	�h[kL�n�yq�n����_e�� -���{H�m��G����}�qw�A��&Z���D�ʞ �aY�SLX�;L��J�ϮN�ZV��)&թ<8�
e�t��|!#���EZ+vq��!�ˤm�{Qb�HL�f�ŘԿir�.�5���J0b��eur��^����3Z�� ���Aɟ��'r�a�/���!��n7�}�	��z�K����n^>��!��(����� �Q�\z�S�T��N��՟x�g�1��oo�����{��Z�+��4_V�H6�o�Tg�#2)�xf�ivѤ|>W�G�"��CN�T6�W<G��I�e��&m4�ޘ|���+;{P������yr̨N��=Q�j�x7Ú�R3e�'Ly��Q��cy�|����
�'��^W�|�}��w�X�=1�`�%(0�ڃ�]^��7#������v�z��3E��RU���iy�؛�4��Ma��G�<zܹ%3b�,|cum�k�C;c8��t.񖳪��?�+%X8��+���J������Y��F>�i�/��D7x��>�Ķ*Kɠ2�D�&���c���>���pe�r&C� ,��Y@����8.4@9A���WH{*�J��]@X+jkeZ6[���f(���s��fSw�h��AL����%�qt�� [���F�7[ΒE�{X��i@������x�(z�wn���;9� �TV<:{�Y�͈�p84u/�F���� '��^OM�1];��g
���:_�"��k@�,�BO)��x{��k���ۼB�N�V��0ZjstsK�Ny�e�?,����y���R�5
 ��t@Vj�f�6����5C�c���t��ʜ
\��d� {�P�v5ޜ'~��c�+I��jy�p�����`�$�-�yl/�zP��p�z(ҧ*����y��k^|�Z0\P���Ɨ�.ʣ}LI�y��>�R�{� �Y��!���O���#�lϸ[�IfnR�M���j�Z�Q�3HM5���]����G��4~���TaҀ��r_���Pٌ�����Xm��6n�0L��?~����T[���9����^ItQ��@idj�Q8E��J���09��?){�a��0�ӄ��f\z��_�'@����n��\��b�|E�\�)�P��-?��Pv�w�� ֫r�6�G��=0�{'����^Hs�gF���mK�0�[L�{�v쒞W�8���.�}ͥ��zv�F:��n���B1��鼇���P�"0n n<�e=蜜����7���ӫ���d.��1m�;����g�+o�����a��˩Ϣ%v�*~�f	}v�d }��RK��#��sB�p�FP�"�}�K�s�,|+�C�2�7�<���9����LR��X����]p�dS0��KM�<�c�>j�,b�E珏:>��#ɨ-[�Q�gʞ�����GEj�[�ƄՍ9 'o!U����/e�]��}i�4���P�e�v_�/~��*nΤn��hrHʜ|0N
��ҧ#�ӣ/�Y+8�Ȉ
�������j^70��.�Y-����Y(��6�D���I�0�Ҿ'ӵ��g���5`���S��&�3p"! DQߣ���cH_2��8}ep^�F�R���k����&,�5P���$������|�I 5�e�vXsHC�ky�t�,F�X����5�3J�ڍU���m)�������v�y���,C�/?
�ohxn}�obUu�I�?\P�$���!Kb���S��XVK>�M�E����B$B�9�#�rN�[7�iq�5Vج�=�@��b2��/�����ظ�����cң'b	_��YwD}c9T�H�)��F��-.�.�]#�\�9
|�T�)nɦ��ӭ3)'�ΥF�O�}Xsd��V`N˃�q�����r2���$!ȪW�v����S���K{�g��{	C>L�%C���7I�i.��m�O� [�����㳔��Zi�@\�`	źXa���c���D	x���NRgvo��*��3K�!T�.m�l�i���"��ZZ�P�GB�U��0�Q���f����W�k��8��[qzR0�~iQւ�>#'m˔�i�>J��uu�5Ʌ@Tt����LA���	,�]���5��F�&9���Έ؟?+He��m9�唨r{qʮ��@HX�2�ܞ$;C*Du�	�p�mU3\h�Ewgx	`����1O����n�CQ�v˲q� �^�}�!ٺI��*�Էq�9uf��R��;�N�Xm��k +:���-��G�^�twnP�Y�/����]u��)jK���1���c&�?pM�*A���'~HTx�k�@�b`r�tY���H��ܘ�`�@�PTT;�ݤ�g����c-r�]�AX'�P�����U ߗ>n}�y`܅����?��#gK9�J����#w�7�����t�R�Li��QAj�"�� Z�t	#'+���;�f�h��Ԧ���
��P��Z���K�
�]͚9�rE$#�|�y;�U���4> iY�-%�g{'��Z��k�qs?�kkg3�zCO�PuNҕO��n�#/�M��[���c<��o�X��Γ��
���th01��9�i����r+h�'�1)�W<p�A)�q��t�~璘:-��� PP���F/�/�T��W	!�i�Z�N�/:L�$��-�ޅ���+�������ڶ���aI�F�<
�
v�C$V>���D�Z �q�Wt�1G��8Y��'®����=��\��rf<�&��;��	km�C7 W������I���4c��\�u��)�{f������[;���c<3���y%���n�W^��ϣb��-�T�+��NQ	^R+����@�Ll����C%�>�ň�e�G�GT��0�]�+��:9?� V?vվߖsS�*�U6t?����z"w~E���ެ�~�	�~/��q�]�ev��Բc5��zZ��X���Reͣ�V� ����cd&=�;����,���c�>< Q2�씮�o-s��H�5�'�~]�ء�d��}<�=�X�G�9s�S�r�,~_���a�H	ۥ��2�&�*w�)�*E?�C��\~�x�e��p488��d�{�&c��5>���FB��#sÆX�=���x�$a򻣰}�-�F�����̨��)��N����z�!sǩ���/�t��[�O螦���i�`s��4�gOg�����-iIk�d3>���'����&eJ}M&9�lsF��d�Xؚ���S �50M&aB��^��6���4x�%$�qA�w�d�O����Ǻ+�vU�B����a������K��NOt曫�^F�S���sD�<��T`���C.[ Ѻ)dN4�6�2�Bz�ݳ�4d.V��v������F��[xS�)&��:�y�G�cb
� /��w�?z��
�ǝ��9�UL�3������#���N���vE�r��P���`	P㛪���PN������i)��@A���ߍ�cmΗ��s���: �DA�EL[�+d �&d6>�5=9���`n0x���s	��l�$a쫦������o�(��>%���4�	x��J�;�+����0(?kB� I]��X�N�0<(�4X�{��xGE��#���]dU����/�/�d�.�L�[�Cqx��e�h��!r�^TB]��X������W��>�2��z��j��ďE�P�="��	N�e^�3A�=�,���8ӱ��lj+�1����Ԡ�}�24[��	�n�=o6�9�Z ��}@\�o�sV��~ @�qٯ�o�ҝ�D��>A)O��/&�¡S���4��G�&�����}P��"������:��~�yl�?�y`BG5 ����=�ߪ��������/����u	.�Oi]N2kx�6���pllT��SF���w�+?n0ܚY5��0l0-����%�̅�qz��������W���n�L�1�^��T�V���_$�=�?b�aֱ�u���?-R����.ɪyG�6�&�=�y~뀕�?؝v4��� dJ�M�O��A�r�����_E��Ed��I!FBBDI�#�.U���],��w���_΢Rp�����`~"��h��V<?G׮�����_�EژW�e�"k=��U
���ëT5��Ÿ�C�R%`����o|\��q�S�'VO�΄���Y����k���0X`Zk�_���oz��&�� ��)���.��㟇~3�>j%��Ot
G�;�ᯜW{�Pk*'����|���o�vi���d�V2��5�i`�!�DY���_��VJz]NR)0�yw�-��3{�;���~/�N,��B�:���A&<�X�I�=AT��V�� �:���hJ:���?���0LE9�b>)�)��[�݋��b\���NDf;���G�B�gȬDh���-�~�3��JW������I�Z�<�f�0���)��3�KE�A�ԄBj��o���]�|�o�/�`&=�K�y���B���#.;~�,`m�4��r�>l5�/�X��������:Zd%��XLt�*�h�0�E?rF)�Kn���R��m�,_A o�O�M�RAi}�����q�����m�)���:�cK���t�y&�O�6(���o��W�\%��x�)M��1pC$6�2�vu��8�ò0M.��F+۸/&l���k8���P�y����~�������䍽~Z[�66	�MX�0�8��}֫�]���ۿ������b~ޤ��8cBXB#d�y�TR�z�i�Iƿ�ت L��Zl�gϺ0l��Ğ?�2�O���a2f�~��)�ÚDT���*p��=� �ّ�z����#jFG����=��7�V���J�v�ed*����ݲ�f#O8d�w[��SS-970>�P��%߇ �n������Ӈ�S4�)f����q��&��&���	F��cH<xG��n?X_�$��� 1 ��ЛCj��^�t��q���#c�O�u�M�"l�
e���t)���BV�d���7x�-�\�x�����(9��t��N�M�5\4�dy�N���LM$5���K>���X|Ճv�X|�?���
`���j��v[�ǻ��D�,t'���6���Jũ�q�lFM ȣg�rI��<�9��w��1MZ��Dd�z�*;:D.���Y�oj��*I��u"���]���I�Ьo�#p���5�;yfnJm������VV�<�&D�$�^�u묮 �S��� ���0K5��(�	�w*S5y�����qW�,w��1�O��4����*�S�$[-(��ڝ�7:�a��o[R��.�Q8����Kݰ��C7|ƴu�l�2}��̅.��/��9"rɉ­[�����w�k.�ڟe7 �z����̋:��m� �8L�/�U�g��a�b"n�۳�������#�7�p��Mca&��8޹��UK��= u� Ƿ׈#x���s%�yqR���65��"���]�ο�ߞ�u�W}na>���ꈚ����l&���t��*�p�t��{p!ziz�a��[O.�p
� ��t9�^�D�̐Ã,��0ts����m�j�C�͹�RΠDPz��lT��:�d�?��Zz�����m��9�4�ج��5Ɔ���������0Sᭋ���mg�@#���Ix/�5F:�ʷ��^2��F��c�J\BYk�|�+.Z0�+��b)�i�2�Ь��~@���ꇨ�*���:�H�/U�m�MUpu�G��xrO�_F����&�m������$���r��w��S_��Ո��W���
��-�YJu��t,!u��J���,�����B�����5�opV�����@x��x��2k�/I��ʝ�iYv}]���	j5�i9ڬΚ]r�4!p�G��=���h��s����(x{�;N}ݮ�;�� p�#��`�	��ZqBL%�0��je�UH��ԑ���L`z)�RHߍk��ʠ��f6�	��iD,��t��vjʵ5��%l�/F��*\M�A��:P.A�n��dDp�s����d�rJa��xX*\������f�ۯ�k��(}�".��ɬ�{r���"<CP[
������Й�ע�{��*���gQ��R�˙�-�cT�����m$������6{�K�	ي1�ﰵ� 4��1�n����{�{q��)��֯5�t�Ct������s�16U�`�t=9#��i$�I�s��^MU�tqOg0l�%r�Ƿd��ߥȀ��0D�Z�B�/���$*=͜���OE��o�0�-�������[@	=��b���s��;�h-�k1�$$�����Ma^�Q��?�*�@�@�:��E	�T�)�4�'��`��:9C���Ԉ���	LvQ�%�����de!Βz���
V����]�pm�^����
	�,}"�ިF���QF~�u#���T����n���d?��>���yz:��TOg��̝�=�d�"�6�$���$�9����<�ȥ������0G�BaY���e����D`uB�*2�1O��� �a���c0㐵�����o�ኵ�KVp4Ԍ��U�A��N���Y�Zm(&%�#��I��Lnz�-�fʶZ��G^����`�oZH�)6zP'1Q̲�n2�d`ş�?� 
v�U�E�����r8�XlxV64EB    cec0    2480���^�ԎX��U�{#c���&���,O"����U[��G�\ki���i^1V��3�H�A�n���c��%�����#r�����P<e�z*��3���q[�&�Jꋻ�~9�V\b���n_T�&�����-)������W�ue�p���FB���DFW�Z��+��.$g"�j.�������* =r� :�6{���E ��(ZB��E��E�{u�f(w��ٳzv]���.?����_2M��u���^�h��x]��}�>43���?�������!7�����%m��u��Hy��+Q�xE��#����wC�L3:%��%�(��h'T�@�T�L�����y#m���U���5�,����w2��&�G������n��׳���!c���Kh��bN�b���$e ��M���_J*�4qI<(����^p����5��x���Ȼ$c��KspřSFIIQ���F��j�)�)z�L?^�V}z{�!��g0����1Ϛ�����҃���$ci�3�\�Qr3�����������;�������]�4@�TRk�̰ �b��"��ő���؃([w�`�� /�&�R6��T���[��7ޮ�n��L�7LՁ�����^��K��-��2|( w�> E9~ݳ/^#TE�we����Nq��� ��I�Ai�>^}�V#)>A���PT5�	,�����3�wb��ӎ��a���)���uoUrF�n�F��{j�k�i:j�V�ě���2�5aGF�]�.O�H.�}��To�І�t�Z��Ͻ[y����D6��%�w��L՘��ʭZ�7,�UY���^�߹T
�D��,(S�GX��W.Y���K
�����2��3��j�F�u�JƗu�R��3���0�8�0�n���Ił*��!��f�G��JB�4��d,sC؇�_l���= �P�T���J��-	�
Ì����S��R��6�P��f�bvT�T� [��kn�Vu���INi���u��t���	������yo^cև3�'�==�����)�gӿ�a�wRH�oQFY ���WM�⿙��[�}�Macl�h��R�5
��{��#�M��]O�-|%?�I��u�L�~�-���$e�T��E������]��Q8ѻna��w0s�b��ȺSBw(�[�{�=�Wβ��S��+7� �z����qH���L"#Ky`p���C�OɊ	� ��ӑX�O.
���I]R~��X�ɲ��I����]<Lɥ64q����}�#>V/��Z�<�+�X�P2�r7!M��Ė��bBdV�̣�gm�A�͔+��Ӛ1jb_Qͧ>d;�h�������#���RfK���3I8��._�d����ɷ���umA�7կ&�+Y�鶔�[��-�
q�����U]��E�RM`0�n�L�ŐV�2 ��.��/���p<j��sۡ\��b��4���6��t�"�g@[Lk��A��~��;����E�m�h}:n؃	����jU�X�� }k[Bf�;S޷l�L-A�?��G�
v��m�Vٞ��K�	���å��M;��C*�
�t4�Q���}ɱ7�~'�B�g���ZH� s��(�b�)�������*�]�P�=]%�{����e�����Y��ᶅj� u�b���e}n/�M�gn�e��c/z����K�8��<_ЪՃ6�m�5Gz�?� �_�-�
5��Z�|���Qd�H�c�k/�=b���ɹ6[�CJ�E(��q���^�ա���4m��؇8q���(x�'Lb��N8�����*�C���2�xO��������Rv_{"��w5��W�_����6�60�����H_�G�|�jd�d�� 
FQް�}��;ג�a������4���ڬ�|���"�|G�R�& x}f'��i�5�'9OI ˏXw�-�{���=$��m}R~� D�h�ըa�k�2�V��K���P�jq��RAm����E�ͫ̄5Q��`E፣\D%J��LX�1ak�S5`U�S�Z�]�D��lI%��)U�kEfk�H����Y���HKP>�R�e��� ��V�P�dd�Hۮ�RV���	Y�����ϔ2mBϏ�f�/������'������^���S��-@N����T�nHخ��e�f����R�@��M�j�_��~l��Qr�&���aD�D2ü"�^�؞�eB(�jH�D�w�㔀��1�`���P���{�	g����x��v��˯�%t.�g�#�C灰���eiG<��DnX�d8��r�=>p��?�}��4�h��5$dY��`�.�V%��p���H�H�}�����~���*�����xK���)�e)f,��4I�X���s��'Y"@����c��cm֜W���� �9�-�<2�n��fo�*���D�*gk�S���>�
[�g�i����8%^�؊.������v���|Q~qxY���m<I��S����݃��X�%] �� �0ܳ�["�`jE'��!R�lͺ���=ߒ�<�DB:��{�e_Ɉ�n��[U�1�pB����`�霘�\@�f��~��L-r�aKrXY��b�q'<M1I�G�=�wWr��+SP�<#ȉ�RhÜ���E�yaVxs�v,Us���p�d֕P=�.R�PY&j�-��:`�����Z��"�-������H�L�S��z��?n�/�l|��Ö>�0�J�b��P!+B"�D��Wt9oki0D�;���HE���J�V'	��W���ox���͐��>�6/[$w�A�enԁ��2�61�w���� ͙�ᾈ��=_�%�3W�12�32��	�G5�0Le����(Hg��L1`Q�cQ��{�4���?�W�<BJF�0���Z�K� d̓�]��{x�����}y2i��
 ���ݵ|m���`��ۂ��,xm��ö�y��#O����q�Ӧ+�ʹU�e�+"���ut�f�<z���"v�ko#"�0(�7#~�d��������Gd3S�#����Cj��>���#b�vGy5Cc�5�uP{�v��������n�����&���"���Td0�l�1�E����1lJ� �A;�LԳ䱼�ٳ�#� y%����,�ey��bPI�t���S0�_.���O��5'��
{�h��`{V:4f�,�P�<_T�1\�!a ���Չ�� dp}�03���o�����h# |��B��aa6%� M�h�=ݙ�>�� ��N4����M% {����s��b�J���_ⳛy���mӸX9�ZY�S�K�!���ݞ�"l���}�$���SG�BA��V���٭����O�əvb ה4=��ه���{ ���p��<�J�5�9��ãߚc�A�b�j:�}�Ƚ $���'�
�����>���#����\�נ"���֋~���`�*�yp�U��H� }L�e0�����%y�G^YM����%WO��l�����ga�}]�d@"z8�1)#�_�U�0��"���d��Q���k�(����jM��l�����"�,HM���x��rr�36*���d|���؁��ĭ�'��PF)�-���Ms��,� ���a� �}��-�\��b�qN'4�H�ls�5�!rS�q���m�AHS�����LA�6Ɍx�2�󰟦�iMR7�I�2��� 6 >���Zb�Պ�lr��������W�թ�
r�n������M���F�Z����Dŧm"}q����17ӥ-���E߮�e���ًw�1g:�Ӟ������N�a�0��e�	���I�c��g9�[�0u|H$b��@�58o�x�~�J�sN�<Z5N:Nl��<�q������3+c�+�:�?3Ø+N���!�J����Yc���T�7����פAEU����c��I�4h�g(y���@B�����]n���8jw)T�'d�a�Ӫɖ�ZW��հ��}%���"fr�����Dxh��E�d�E��y�C֮~�:�Bc*oQ��r�`Ą猉�H|��8�-'�*�k�{���-]^�t�f&"w��SmD{gt%��LmX�(��q��N���WO��R�%+��7�6?n�X;Bzm.>c�C�4�ޙ��m�$�T�ǚF��o����J�@Ӝz�]J���=7E>C>6��nA۵�d�A��`��O�㍷��;9���_S��r4�A,��G=p�27����ڌ��p������x������
e���o���U��2�/�E{�|v]������޷�c�*��{�T��L	�z�����D���W���s�՝�A�����m�o�~K7�Z� �w ��0����{�6�D݄˰��[�zܐ6l����\��<F�O���܏�/Q�>&qLUoTvÐ�q �?s���4^�m5޻Vp��Ҹ�/�c�1�O�+
Ί�.�lf׿��OL@�E1�'����_��7�9�QQ�����͌��b8H�C��)����v���}�����:���^�*����}�z��{sa�Y#�$|�ɫ�Zp�^��`B45Ƭ`����}g9���#}k��C�[;�V`��_�No�ʏ�*�(�7���ŏ��ws�r�!���؝�KH��U���mR,�+�<w��:e��E{f����A���7�7w�a�<�KL��YKt������	����P�-�8�.ٌcb*u�ѯ�=�-|ʖ'�RO���=��f���������.�y?�'l(��=�(,�G�V���^?�q��ޓ<����u�X�Ҋ5~�X���4I,���Gi+<ꄶK�.Z^�0ƫ��rz\����,:qR�ǅ���K�#���܌�6�٫0��w����
ո�!�N*�aVuU8�����<%"��k."�!-y���G.�L���ª��d5����ٶ��sPb�~Ǜɦu�t+���Uz�V��(q�Z�c�'�C�<���@�VA�u�����~���h�%�Ը}��a~n]�G(-�E�V(����)
H)�[�
w����� ![wb��>��@EtR/y5�HP>x����6�����Fw����|��wQ����<�/�a��|��Ǯc��k��D�Skޜ�1&��?�B-�{yU�N�2�"FDna��wz��̺:�O�-@v��E_�v&'z��R*rf J���b  "m����]�_�ȷ�J�pa�}X>/���u�c�w,�����wC;J}X�1V0��y-zjOz��Y;�}P+� ����>�c2�	~%����FpP�X$�����<��]K�g���;g����T�Q���񾅙����k�[wJ�|�[a�C՜B�o��e;���1�ެ�J@f��R
|-j��E}��q�1�I������fm���[?m�Q��6������R]U��퍵�Uղ�?�U���후���0��ҥX\��۩�!qn����z���8;�F�#�0S�[c΄�RV�'\ֲN{ݮ�w�А�&�aZ�a�)��	c,��X���G����淽��7ψ�ܩV�\��#D�I�Խ��&i��*��S�Ϣ�v4��%o8BLqy�n�6�}E���=�p-d�Х�0�vK��Zd}}�#w�B��o1�bW�R�iC�VEI;��hi�+�:P����Y$�=	项V��P$x���r}�i4?���g��=�)�o?�X<�V�Z�����7�*��VqK�i:�ݧf����.u`���r_l�/�q|샙�aa��/*����S������U8��!����0hd���s5��K���M��D���;������Gy$қ��h�W�(ӡ�p�w�=*�36�մd�C�,y�{9Fx�4���z�Y�"��Z���u[�W��]d$�6D�壆k��=�+z�H?C��I�jSȩPj��y��-�����*��.s���tE��iG�w>���������E!�ϒ3<��e�W�*|�R��e�
��'Lm ��#)$�w����)v'�M������_%�� e�0��76P��0����)H��_����x�kJf`6l��XD�'���a1��S�RLM�C��l0�&��k%��I}q�������?���*��P�D�@ַQ�G��2S��ch�X�AG5��eM�����G�����(Ni��f�s�U�	Z�ڔ�nB)3�HȮ��Az�������&��/����{#�R9�.�9N`}�4�}��3`F�i������6��ʒ�o<�1~$e����y�@�(@� �?J�[f��:�7��F^������7�8~���Dk.7�0�F�+i����+dq{>@�hQ��x%�9*����i[F����U�+�e��G��Cw���Ni-Y���Py1G2�=cɘ(t���}%/��g�I�9pA%��uc��gc�+=ٲC���;��c�o�RQ��,ة���c��<rLwG �i�;��ސP�P�J�(��p�@A﫞���H�C-�qRd��Ot�E�[`!F]
�.���hd�E,/���ˀ��F�%�T�	|>����!{�n�k/S���vMYj^�?O�sMv�#�!��
��������w4Dg�8���T�������kɼ��|�وl�.ף�O�"%6YֿTv4���q�s'���8�e�1T��\!ˎ��џ��J�d�]��rn�����l�f�Z��|���
pa�H����;aA�^�Z ���~����}O�Ɖp�rU�P3��:�L�8�*pV4���r!�{sI�ܾ��ōB��,P����� �θ��jq[��_����ԎoJ8�=^�f�EY��4�5(��l�����f��r5�N� ~���U:;�;�C�~���/����W�̟&v�Ò�-M7���U�ۑo����l���8���@ҳ�M�5�����|6:�j;����#�X�x�?�%9��n�7�g#���;}�;Ѐ���va���FھRZ:�Z��.@a�f�@���޴{m�њќW���Z;U�O� *\KR���l��ݒN�<7��n���>��zPJs�\�J�;����O�(4����s���S�#g��
�e&�-����@'�"r�r4�-2!u;QA�ڱ~OO��z&�P��"�l�ro�|V����b��������G�B�^?��|��Lu6�� �/b6��+�6*b�K���\�G�����5��Ѽ��8�]��;���ͼ	��W�/O�U�?pS���V�P��H�O���c����	�gg�A[�K��6י-��m^�Y �����LKJqF0��V��E���]������e=�����Un�_ׯ��@C�G�f�ĖЛ�	��Z�c45��9�z��ѧ�)i<�?��5X�,��X>G&e�S�@,��R��א�~�epJw�����{kV:�!Ʃ'!t�GL��wx�o�^/�B<�8Ӄpj �`�M��Ϗ�cS���k�g낌�5��C��}�U�����?!;��֜�N��Ud�9�y�~�� �[�RZ�
SB�����F���n"9���u�e<�Ș�P�"�:�y��P�՗��|K=�%�[�e% 3�έf�v����{ө̡h�=T<@
����q�mK��|�rTE��RF�p�ѕ�`?2������q�;���V���=k��s�N
�̨+L�æʝB0+k��%��e���T]M�~c \r��u��ַ��3�?���i�����O'�!<��/:9�'��ܐ�<S�����y/�Ԗm��13M�:�D\�
���$6r1��|�{�e�-��F��ꥇ���X"q)y@^r_*��Zִ�7��ՠ[e�:��^i�����T4�}
�r {nz4*÷׆�z���$�Q��(Z�U�\�h0�̴ �7<o��҃H�ܞ��Y�p �(���h��=�7z����.�=�kHie�DZ��ʊ>�Ǘ��d�>Q�(1DG������uT4�������� *�����XO�ǰk�低�ţ9��ң1(o�RA�(�M�S	9�����r�7X�f�;\A+<�XH�<l'z�,�K�lDiM;��+��UnX�x͋-��V�(���P�nzs���03�=U��EkS�&�-!vK��b�B��|*�3��yMY2�&ޙ���c@znƝ�� �;.�YI��=�a�~~���]��i��Y�]#�=���6�^��ןH��>�1��>��t�ڛ�ή��?y������B��i9e�t�Bΐj��~�a�Qx�<�-!�:�-����c�C�n�&i 6O���u\U� ��knJ�'���w�yFC�:��''��?v���.�H\�o:�)��KW��uD��d�M�/Q�X .	&��ǆ.��Ȅ��E�t<�X�RH����M;1kf���+��E��-O�Z`L<J�e:u�X�mv�Z1�\3m��V"�{�D�}4��'<�Q�K��O3~qu)FB���b�g�Ir��ڂ��?v;v'�*���G��f�\����ZW��OU�<)��s�T1�~$�MT,|��Y�w4�T����z;4Ш�1���'9��?�긐�W�4sIv���\�ߕ���A �T��m��̨�J�ɞP�S:��!*��1�@�RF>��n��j���m�z'}<�HTfg5ٸ{��M���_��!��y��B �����r��?���pd�'E��z/�%td/�㸋�eC}���ah~9�8�C��X��q���:��S������l�2o�_8啣~����oB�HQB��J@E��h1gp�و�`؏m̌�@k����6�y�B�}F�᫓���ۋ���w8U<����� ��̄�˜�˗Ÿ�q�S���g��Kљ��c1���40GE���A���\����rq/�2 ��!�rAU�C����-u�@���U�d�<ɭ�;M����_��� 2��s5J���?'Fx��PaK?��{!��f��Б�xp�3���[������fak�ꣾ��k���\̩̲3�F�T�b#m��)�v+�B��jn|�y?�1H��O��T�;&5̐+�V��r�O-��,��<(g��~���k)���2���t����*�h�j�I����Y����� _=�)5N�������܂]�k��$�p�d)m�L��!<U��抷���!M�>s��LOf�tY�����5�� =�������B�3�<;���>zC���,%����Yg����*k�y.��