XlxV64EB    1595     840�z6=.~t���P���t�c��l׀vO��5����P�㉻�a5|�6o��:�^$��>��	EB��[g��� *��-rd ����~>��/��s:l���۫��4�'G����0�X����omr��,�bZCߏ����4� pG� 6C^p y`��<
p�~i���5���St���G�26`p�g{����?ۆ���e��S&/C�A��)Y�u^F���L���=�^?�l��J�<cg̋���ٱD��V1jHm����Zٹ����w���L����-DR�'�@.R�~Ķ-@,�`0�Q��S��9����v�6���^YA0>����fO~��Bn����S데��m�mW*�	Hܸ��O�=M��������f*��F4!�W
U�u꽟|1�����}�J �@���K�*���<����T��WgњS�c��"�~�2t��p�D8� '�&�#���/UΦv�X���
���@N�T�b�;5�^���7�\����~]�����of����Q��2-U�+_��IY�����87����f+Sڇ-q��\�4Z�-] Ce9l�h�e;u�F��j��i\���y��Q:@�ϋ4�Ư�z�l�4����ԌXc���f�2r&�j�U�����q�?�=Ҙ�,�h�yq5��h>�Z����~Ұg�p�TBw���Aad�ګ�q�`w�h}|N��N��}ّ.����������[�t�/�����'�N�ƯP�y��KX0��w��_�����g}ǝ�|s�'�A�H�q���M3�vF.�&I��TT�_Km�yz�"�)"��{���\=J�i�6T�`y9A*�i3���!��_*T����.�u�#v~mO�.l�� �&��&M�m�
?N�0�DO�3�D]�-�ԉx��]���3ukwJ�"q��TX
��ɯ=ܫ�>^���_�x�H\���>{�R4 �u'̓dPV"
���N͢oK�m�Ph/|�0�%�=�Z��Op���"�p����]ܶ&�Jd7~pC�x�~�EIo�	l��3C��(c(4l7a�3|("���}LR%�,op ���i"��`K\(�e	Tl�H!�ݮt
_
�tR�M���<�c�3!D�Z�����WȆEi�@�?s$�n-��Si������E�l��A��iU�F�r5���l����먺��7�3�o���<����~��4]j	D�A�,�z�ܱ!f0�� �N,�@�[;�d�N� �Ղ�]2��ӦRL�i���2�ޅ���~�����D�V8���GI�����N~����y���p��WH�=�4���֑���oo���M�C/�Czl���g��A��:�2���:��c�JTw�A�Y|P�݊#7��\,�_�Jx�S�]��������3�&iv�dQ1J,hZ�z��Ma�k���p��_샹����=!
�GK2�F">�g��ϰb�Y�����Οd�v�2!lK��$�� ���N��}�|U�X�FkP�9/�`]G1�	N����mǯD�v�XȮ�әĔoK��~�5JSv�#,������*��j�����eG|imq%�H�����<sp8޲8�W���(Y�<�v�kL�V��8v�r���Sl���0
^u�x�Ww�~�
'�z^|E�b��g^ �1�Z+S��
�U`n� &�%�C��<-9\Ҽ� T��1]�qD����2�1��O� N��#�u��^O�VN�n�X=�V�^�8H^�J%~����;'�SG����(�	�#3�[lŮO�Xd��F�W��ϥb3h�ZA��0�#����H$�N��f���sNg�"9].�]�������׽��:��gwE^��ឣK�ŒY�=�b���c$���pXf�_p��]�}�q�[Y�@���e������L�yM��J@�\���kּcf�岥�m�����C��5���U��E�0�9?~0���ƮU���=���ϯ$�zժ�z�%M��Y�%��ҳ��cbl��Ʉ�KU觘��?R��p�b��#�J���Fڴ2,h������C�%�k��J]J���!O�/�